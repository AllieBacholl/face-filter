module immediate_execution(

    input [24:0] instruction_without_opcode,
    input [2:0] imm_ctrl_ID,
    output logic [31:0] imm_res_ID
);



endmodule
