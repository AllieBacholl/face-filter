module systolic_controller
#(

)
(
    input done,
    output clr,
    output start,

);
endmodule