module immediate_execution(

    input logic [24:0] instruction_wo_opcode,
);



endmodule
