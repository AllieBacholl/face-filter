module UART_control (
    input clk,
    input rst_n,
    input tbr,
    input rx_
)