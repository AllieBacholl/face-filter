module tb_img2col8();
    
endmodule