// bram.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module bram (
		input  wire        clk_clk,               //        clk.clk
		input  wire [9:0]  mem_data_0_address,    // mem_data_0.address
		input  wire        mem_data_0_clken,      //           .clken
		input  wire        mem_data_0_chipselect, //           .chipselect
		input  wire        mem_data_0_write,      //           .write
		output wire [63:0] mem_data_0_readdata,   //           .readdata
		input  wire [63:0] mem_data_0_writedata,  //           .writedata
		input  wire [7:0]  mem_data_0_byteenable, //           .byteenable
		input  wire [9:0]  mem_data_1_address,    // mem_data_1.address
		input  wire        mem_data_1_chipselect, //           .chipselect
		input  wire        mem_data_1_clken,      //           .clken
		input  wire        mem_data_1_write,      //           .write
		output wire [63:0] mem_data_1_readdata,   //           .readdata
		input  wire [63:0] mem_data_1_writedata,  //           .writedata
		input  wire [7:0]  mem_data_1_byteenable, //           .byteenable
		input  wire [9:0]  mem_data_2_address,    // mem_data_2.address
		input  wire        mem_data_2_clken,      //           .clken
		input  wire        mem_data_2_chipselect, //           .chipselect
		input  wire        mem_data_2_write,      //           .write
		output wire [63:0] mem_data_2_readdata,   //           .readdata
		input  wire [63:0] mem_data_2_writedata,  //           .writedata
		input  wire [7:0]  mem_data_2_byteenable, //           .byteenable
		input  wire [9:0]  mem_data_3_address,    // mem_data_3.address
		input  wire        mem_data_3_chipselect, //           .chipselect
		input  wire        mem_data_3_clken,      //           .clken
		input  wire        mem_data_3_write,      //           .write
		output wire [63:0] mem_data_3_readdata,   //           .readdata
		input  wire [63:0] mem_data_3_writedata,  //           .writedata
		input  wire [7:0]  mem_data_3_byteenable, //           .byteenable
		input  wire        reset_reset_n          //      reset.reset_n
	);

	wire    rst_controller_reset_out_reset;     // rst_controller:reset_out -> [onchip_memory2_0:reset, onchip_memory2_0:reset2, onchip_memory2_1:reset, onchip_memory2_1:reset2]
	wire    rst_controller_reset_out_reset_req; // rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, onchip_memory2_1:reset_req, onchip_memory2_1:reset_req2]

	bram_onchip_memory2_0 onchip_memory2_0 (
		.clk         (clk_clk),                            //   clk1.clk
		.address     (mem_data_0_address),                 //     s1.address
		.clken       (mem_data_0_clken),                   //       .clken
		.chipselect  (mem_data_0_chipselect),              //       .chipselect
		.write       (mem_data_0_write),                   //       .write
		.readdata    (mem_data_0_readdata),                //       .readdata
		.writedata   (mem_data_0_writedata),               //       .writedata
		.byteenable  (mem_data_0_byteenable),              //       .byteenable
		.reset       (rst_controller_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req), //       .reset_req
		.address2    (mem_data_1_address),                 //     s2.address
		.chipselect2 (mem_data_1_chipselect),              //       .chipselect
		.clken2      (mem_data_1_clken),                   //       .clken
		.write2      (mem_data_1_write),                   //       .write
		.readdata2   (mem_data_1_readdata),                //       .readdata
		.writedata2  (mem_data_1_writedata),               //       .writedata
		.byteenable2 (mem_data_1_byteenable),              //       .byteenable
		.clk2        (clk_clk),                            //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                // (terminated)
	);

	bram_onchip_memory2_1 onchip_memory2_1 (
		.clk         (clk_clk),                            //   clk1.clk
		.address     (mem_data_2_address),                 //     s1.address
		.clken       (mem_data_2_clken),                   //       .clken
		.chipselect  (mem_data_2_chipselect),              //       .chipselect
		.write       (mem_data_2_write),                   //       .write
		.readdata    (mem_data_2_readdata),                //       .readdata
		.writedata   (mem_data_2_writedata),               //       .writedata
		.byteenable  (mem_data_2_byteenable),              //       .byteenable
		.reset       (rst_controller_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req), //       .reset_req
		.address2    (mem_data_3_address),                 //     s2.address
		.chipselect2 (mem_data_3_chipselect),              //       .chipselect
		.clken2      (mem_data_3_clken),                   //       .clken
		.write2      (mem_data_3_write),                   //       .write
		.readdata2   (mem_data_3_readdata),                //       .readdata
		.writedata2  (mem_data_3_writedata),               //       .writedata
		.byteenable2 (mem_data_3_byteenable),              //       .byteenable
		.clk2        (clk_clk),                            //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
