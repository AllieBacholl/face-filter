module interrupt_handler(
    input clk, rst,
    input external,
    output interrupt_handling_addr,
    output interrupt_ctrl
);
    
endmodule