// https://github.com/AllieBacholl/face-filter.git

module proc(
    input clk, RST, EXT
    output err
);



endmodule