// *****************************************************************************
//
// Copyright 2007-2016 Mentor Graphics Corporation
// All Rights Reserved.
//
// THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE PROPERTY OF
// MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS.
//
// *****************************************************************************
// SystemVerilog           Version: 20160107
// *****************************************************************************

// Title: axi_top
//

package mgc_axi_pkg;
import QUESTA_MVC::*;

`ifdef MODEL_TECH
// *****************************************************************************
//
// Copyright 2007-2016 Mentor Graphics Corporation
// All Rights Reserved.
//
// THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE PROPERTY OF
// MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS.
//
// *****************************************************************************
// SystemVerilog           Version: 20160107
// *****************************************************************************

// Title: AXI Enumeration Types
//

//------------------------------------------------------------------------------
//
// Enum: axi_size_e
//
//------------------------------------------------------------------------------
//  Word size encoding 
typedef enum bit [2:0]
{
    AXI_BYTES_1   = 3'h0,
    AXI_BYTES_2   = 3'h1,
    AXI_BYTES_4   = 3'h2,
    AXI_BYTES_8   = 3'h3,
    AXI_BYTES_16  = 3'h4,
    AXI_BYTES_32  = 3'h5,
    AXI_BYTES_64  = 3'h6,
    AXI_BYTES_128 = 3'h7
} axi_size_e;



//------------------------------------------------------------------------------
//
// Enum: axi_prot_e
//
//------------------------------------------------------------------------------
//  Protection type 
typedef enum bit [2:0]
{
    AXI_NORM_SEC_DATA    = 3'h0,
    AXI_PRIV_SEC_DATA    = 3'h1,
    AXI_NORM_NONSEC_DATA = 3'h2,
    AXI_PRIV_NONSEC_DATA = 3'h3,
    AXI_NORM_SEC_INST    = 3'h4,
    AXI_PRIV_SEC_INST    = 3'h5,
    AXI_NORM_NONSEC_INST = 3'h6,
    AXI_PRIV_NONSEC_INST = 3'h7
} axi_prot_e;



//------------------------------------------------------------------------------
//
// Enum: axi_cache_e
//
//------------------------------------------------------------------------------
//  Cache type
typedef enum bit [3:0]
{
    AXI_NONCACHE_NONBUF             = 4'h0,
    AXI_BUF_ONLY                    = 4'h1,
    AXI_CACHE_NOALLOC               = 4'h2,
    AXI_CACHE_BUF_NOALLOC           = 4'h3,
    AXI_CACHE_RSVD0                 = 4'h4,
    AXI_CACHE_RSVD1                 = 4'h5,
    AXI_CACHE_WTHROUGH_ALLOC_R_ONLY = 4'h6,
    AXI_CACHE_WBACK_ALLOC_R_ONLY    = 4'h7,
    AXI_CACHE_RSVD2                 = 4'h8,
    AXI_CACHE_RSVD3                 = 4'h9,
    AXI_CACHE_WTHROUGH_ALLOC_W_ONLY = 4'ha,
    AXI_CACHE_WBACK_ALLOC_W_ONLY    = 4'hb,
    AXI_CACHE_RSVD4                 = 4'hc,
    AXI_CACHE_RSVD5                 = 4'hd,
    AXI_CACHE_WTHROUGH_ALLOC_RW     = 4'he,
    AXI_CACHE_WBACK_ALLOC_RW        = 4'hf
} axi_cache_e;



//------------------------------------------------------------------------------
//
// Enum: axi_burst_e
//
//------------------------------------------------------------------------------
//  This specifies Burst type which determines address calculation
typedef enum bit [1:0]
{
    AXI_FIXED      = 2'h0,
    AXI_INCR       = 2'h1,
    AXI_WRAP       = 2'h2,
    AXI_BURST_RSVD = 2'h3
} axi_burst_e;



//------------------------------------------------------------------------------
//
// Enum: axi_response_e
//
//------------------------------------------------------------------------------
//  Response type 
typedef enum bit [1:0]
{
    AXI_OKAY   = 2'h0,
    AXI_EXOKAY = 2'h1,
    AXI_SLVERR = 2'h2,
    AXI_DECERR = 2'h3
} axi_response_e;



//------------------------------------------------------------------------------
//
// Enum: axi_lock_e
//
//------------------------------------------------------------------------------
//  Lock type for atomic accesses
typedef enum bit [1:0]
{
    AXI_NORMAL    = 2'h0,
    AXI_EXCLUSIVE = 2'h1,
    AXI_LOCKED    = 2'h2,
    AXI_LOCK_RSVD = 2'h3
} axi_lock_e;



//------------------------------------------------------------------------------
//
// Enum: axi_rw_e
//
//------------------------------------------------------------------------------
//  Specifies transaction type read or write 
typedef enum bit [0:0]
{
    AXI_TRANS_READ  = 1'h0,
    AXI_TRANS_WRITE = 1'h1
} axi_rw_e;



//------------------------------------------------------------------------------
//
// Enum: axi_len_e
//
//------------------------------------------------------------------------------
//  Specifies length of the transaction 
typedef enum bit [3:0]
{
    AXI_LENGTH_1  = 4'h0,
    AXI_LENGTH_2  = 4'h1,
    AXI_LENGTH_3  = 4'h2,
    AXI_LENGTH_4  = 4'h3,
    AXI_LENGTH_5  = 4'h4,
    AXI_LENGTH_6  = 4'h5,
    AXI_LENGTH_7  = 4'h6,
    AXI_LENGTH_8  = 4'h7,
    AXI_LENGTH_9  = 4'h8,
    AXI_LENGTH_10 = 4'h9,
    AXI_LENGTH_11 = 4'ha,
    AXI_LENGTH_12 = 4'hb,
    AXI_LENGTH_13 = 4'hc,
    AXI_LENGTH_14 = 4'hd,
    AXI_LENGTH_15 = 4'he,
    AXI_LENGTH_16 = 4'hf
} axi_len_e;



//------------------------------------------------------------------------------
//
// Enum: axi_error_e
//
//------------------------------------------------------------------------------
//  Specifies error type 
typedef enum bit [3:0]
{
    AXI_AWBURST_RSVD        = 4'h0,
    AXI_ARBURST_RSVD        = 4'h1,
    AXI_AWSIZE_GT_BUS_WIDTH = 4'h2,
    AXI_ARSIZE_GT_BUS_WIDTH = 4'h3,
    AXI_AWLOCK_RSVD         = 4'h4,
    AXI_ARLOCK_RSVD         = 4'h5,
    AXI_AWLEN_LAST_MISMATCH = 4'h6,
    AXI_AWID_WID_MISMATCH   = 4'h7,
    AXI_WSTRB_ILLEGAL       = 4'h8,
    AXI_AWCACHE_RSVD        = 4'h9,
    AXI_ARCACHE_RSVD        = 4'ha
} axi_error_e;



//------------------------------------------------------------------------------
//
// Enum: axi_assertion_e
//
//------------------------------------------------------------------------------
//  Type defining the assertion messages which can be produced by the <mgc_axi> QVIP.
// 
// Individual assertion messages can be disabled using the <config_enable_assertion> array of configuration bits.
// 
// AXI_ARESETn_SIGNAL_Z                                                        -  60000 -  AXI reset signal (ARESETn) has a value Z
// AXI_ARESETn_SIGNAL_X                                                        -  60001 -  AXI reset signal (ARESETn) has a value X
// AXI_ACLK_SIGNAL_Z                                                           -  60002 -  
// AXI_ADDR_FOR_READ_BURST_ACROSS_4K_BOUNDARY                                  -  60004 -  This read transaction has crossed a 4KB boundary (SPEC3(A3.4.1))
// AXI_ADDR_FOR_WRITE_BURST_ACROSS_4K_BOUNDARY                                 -  60005 -  This write transaction has crossed a 4KB boundary (SPEC3(A3.4.1))
// AXI_ARADDR_CHANGED_BEFORE_ARREADY                                           -  60006 -  The value of <ARADDR> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARADDR_UNKN                                                             -  60007 -  <ARADDR> has an X value/<ARADDR> has an Z value (SPEC3(A2.5))
// AXI_ARBURST_CHANGED_BEFORE_ARREADY                                          -  60008 -  The value of <ARBURST> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARBURST_UNKN                                                            -  60009 -  <ARBURST> has an X value/<ARBURST> has an Z value (SPEC3(A2.5))
// AXI_ARCACHE_CHANGED_BEFORE_ARREADY                                          -  60010 -  The value of <ARCACHE> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARCACHE_UNKN                                                            -  60011 -  <ARCACHE> has an X value/<ARCACHE> has an Z value (SPEC3(A2.5))
// AXI_ARID_CHANGED_BEFORE_ARREADY                                             -  60012 -  The value of <ARID> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARID_UNKN                                                               -  60013 -  <ARID> has an X value/<ARID> has an Z value (SPEC3(A2.5))
// AXI_ARLEN_CHANGED_BEFORE_ARREADY                                            -  60014 -  The value of <ARLEN> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARLEN_UNKN                                                              -  60015 -  <ARLEN> has an X value/<ARLEN> has an Z value (SPEC3(A2.5))
// AXI_ARLOCK_CHANGED_BEFORE_ARREADY                                           -  60016 -  The value of <ARLOCK> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARLOCK_UNKN                                                             -  60017 -  <ARLOCK> has an X value/<ARLOCK> has an Z value (SPEC3(A2.5))
// AXI_ARPROT_CHANGED_BEFORE_ARREADY                                           -  60018 -  The value of <ARPROT> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARPROT_UNKN                                                             -  60019 -  <ARPROT> has an X value/<ARPROT> has an Z value (SPEC3(A2.5))
// AXI_ARREADY_UNKN                                                            -  60020 -  <ARREADY> has an X value/<ARREADY> has a Z value (SPEC3(A2.5))
// AXI_ARSIZE_CHANGED_BEFORE_ARREADY                                           -  60021 -  The value of <ARSIZE> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARSIZE_UNKN                                                             -  60022 -  <ARSIZE> has an X value/<ARSIZE> has an Z value (SPEC3(A2.5))
// AXI_ARUSER_CHANGED_BEFORE_ARREADY                                           -  60023 -  The value of <ARUSER> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARUSER_UNKN                                                             -  60024 -  <ARUSER> has an X value/<ARUSER> has an Z value (SPEC3(A2.5))
// AXI_ARVALID_DEASSERTED_BEFORE_ARREADY                                       -  60025 -  <ARVALID> has been de-asserted before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                 -  60026 -  A master interface must begin driving <ARVALID> high only at a rising clock edge after <ARESETn> is HIGH (SPEC3(A3.1.2))
// AXI_ARVALID_UNKN                                                            -  60027 -  <ARVALID> has an X value/<ARVALID> has an Z value (SPEC3(A2.5))
// AXI_AWADDR_CHANGED_BEFORE_AWREADY                                           -  60028 -  The value of <AWADDR> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))
// AXI_AWADDR_UNKN                                                             -  60029 -  <AWADDR> has an X value/<AWADDR> has an Z value (SPEC3(A2.2))
// AXI_AWBURST_CHANGED_BEFORE_AWREADY                                          -  60030 -  The value of <AWBURST> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))
// AXI_AWBURST_UNKN                                                            -  60031 -  <AWBURST> has an X value/<AWBURST> has an Z value (SPEC3(A2.2))
// AXI_AWCACHE_CHANGED_BEFORE_AWREADY                                          -  60032 -  The value of <AWCACHE> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                       
// AXI_AWCACHE_UNKN                                                            -  60033 -  <AWCACHE> has an X value/AWCACHE has an Z value (SPEC3(A2.2))
// AXI_AWID_CHANGED_BEFORE_AWREADY                                             -  60034 -  The value of <AWID> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))
// AXI_AWID_UNKN                                                               -  60035 -  <AWID> has an X value/<AWID> has an Z value (SPEC3(A2.2))
// AXI_AWLEN_CHANGED_BEFORE_AWREADY                                            -  60036 -  The value of <AWLEN> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))
// AXI_AWLEN_UNKN                                                              -  60037 -  <AWLEN> has an X value/<AWLEN> has an Z value (SPEC3(A2.2))                                                                                                                                        
// AXI_AWLOCK_CHANGED_BEFORE_AWREADY                                           -  60038 -  The value of <AWLOCK> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                            
// AXI_AWLOCK_UNKN                                                             -  60039 -  <AWLOCK> has an X value/<AWLOCK> has an Z value (SPEC3(A2.2))
// AXI_AWPROT_CHANGED_BEFORE_AWREADY                                           -  60040 -  The value of <AWPROT> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                          
// AXI_AWPROT_UNKN                                                             -  60041 -  <AWPROT> has an X value/<AWPROT> has an Z value (SPEC3(A2.2))                                                                                                                                        
// AXI_AWREADY_UNKN                                                            -  60042 -  <AWREADY> has an X value/<AWREADY> has an Z value (SPEC3(A2.2))                                                                                                                                        
// AXI_AWSIZE_CHANGED_BEFORE_AWREADY                                           -  60043 -  The value of <AWSIZE> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                                       
// AXI_AWSIZE_UNKN                                                             -  60044 -  <AWSIZE> has an X value/<AWSIZE> has an Z value (SPEC3(A2.2))                                                                                                                                                 
// AXI_AWUSER_CHANGED_BEFORE_AWREADY                                           -  60045 -  The value of <AWUSER> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                                           
// AXI_AWUSER_UNKN                                                             -  60046 -  <AWUSER> has an X value/<AWUSER> has an Z value (SPEC3(A3.1))                                                                                                                                                    
// AXI_AWVALID_DEASSERTED_BEFORE_AWREADY                                       -  60047 -  <AWVALID> has been de-asserted before <AWREADY> was asserted (SPEC3(A3.2.2))                                                                                                                  
// AXI_AWVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                 -  60048 -  A master interface must begin driving <AWVALID> high only at a rising clock edge after <ARESETn> is HIGH (SPEC3(A3.1.2))                                                               
// AXI_AWVALID_UNKN                                                            -  60049 -  <AWVALID> has an X value/<AWVALID> has an Z value (SPEC3(A2.2))                                                                                                                                                 
// AXI_BID_CHANGED_BEFORE_BREADY                                               -  60050 -  The value of <BID> has changed from its initial value between the time <BVALID> was asserted, and before <BREADY> was asserted (SPEC3(A3.2.1))                                                 
// AXI_BID_UNKN                                                                -  60051 -  <BID> has an X value/<BID> has a Z value (SPEC3(A2.4))                                                                                                                                                       
// AXI_BREADY_UNKN                                                             -  60052 -  <BREADY> has an X value/<BREADY> has an Z value (SPEC3(A2.4))                                                                                                                                                 
// AXI_BRESP_CHANGED_BEFORE_BREADY                                             -  60053 -  The value of <BRESP> has changed from its initial value between the time <BVALID> was asserted, and before <BREADY> was asserted (SPEC3(A3.2.1))                                            
// AXI_BRESP_UNKN                                                              -  60054 -  <BRESP> has an X value/<BRESP> has a Z value (SPEC3(A2.4))                                                                                                                                                   
// AXI_BUSER_CHANGED_BEFORE_BREADY                                             -  60055 -  The value of <BUSER> has changed from its initial value between the time <BVALID> was asserted, and before <BREADY> was asserted (SPEC3(A3.2.1))                                       
// AXI_BUSER_UNKN                                                              -  60056 -  <BUSER> has an X value/<BUSER> has a Z value (SPEC3(A2.4))                                                                                                                                                       
// AXI_BVALID_DEASSERTED_BEFORE_BREADY                                         -  60057 -  <BVALID> has been de-asserted before <BREADY> was asserted (SPEC3(A3.2.1))                                                                                                                       
// AXI_BVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  -  60058 -  A slave interface must begin driving  <BVALID> high only at a rising clock edge after ARESETn is HIGH (SPEC3(A3.1.2))                                                                        
// AXI_BVALID_UNKN                                                             -  60059 -  <BVALID> has an X value/<BVALID> has a Z value (SPEC3(A2.4))                                                                                                                                                   
// AXI_EXCLUSIVE_READ_ACCESS_MODIFIABLE                                        -  60060 -  The modifiable bit (bit 1 of the cache parameter) should not be set for an exclusive read access (SPEC3(A7.2.4))                                                                                 
// AXI_EXCLUSIVE_READ_BYTES_TRANSFER_EXCEEDS_128                               -  60061 -  Number of bytes in an exclusive read transaction must be less than or equal to 128 (SPEC3(A7.2.4))                                                                                         
// AXI_EXCLUSIVE_WRITE_BYTES_TRANSFER_EXCEEDS_128                              -  60062 -  Number of bytes in an exclusive write transaction must be less than or equal to 128 (SPEC3(A7.2.4))                                                                                
// AXI_EXCLUSIVE_READ_BYTES_TRANSFER_NOT_POWER_OF_2                            -  60063 -  Number of bytes of an exclusive read transaction is not a power of 2 (SPEC3(A7.2.4))                                                                                           
// AXI_EXCLUSIVE_WRITE_BYTES_TRANSFER_NOT_POWER_OF_2                           -  60064 -  Number of bytes of an exclusive write transaction is not a power of 2 (SPEC3(A7.2.4))                                                                                               
// AXI_EXCLUSIVE_WR_ADDRESS_NOT_SAME_AS_RD                                     -  60065 -  Exclusive write does not match the address of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                                        
// AXI_EXCLUSIVE_WR_BURST_NOT_SAME_AS_RD                                       -  60066 -  Exclusive write does not match the burst setting of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                                      
// AXI_EXCLUSIVE_WR_CACHE_NOT_SAME_AS_RD                                       -  60067 -  Exclusive write does not match the cache setting of the previous exclusive read to this id (see the ARM AXI compliance-checker AXI_RECM_EXCL_MATCH assertion code) (SPEC3(A7.2.4))            
// AXI_EXCLUSIVE_WRITE_ACCESS_MODIFIABLE                                       -  60068 -  The modifiable bit (bit 1 of the cache parameter) should not be set for an exclusive write access (SPEC3(A7.2.4))                                                               
// AXI_EXCLUSIVE_WR_LENGTH_NOT_SAME_AS_RD                                      -  60069 -  Exclusive write does not match the length of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                           
// AXI_EXCLUSIVE_WR_PROT_NOT_SAME_AS_RD                                        -  60070 -  Exclusive write does not match the prot setting of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                       
// AXI_EXCLUSIVE_WR_SIZE_NOT_SAME_AS_RD                                        -  60071 -  Exclusive write does not match the size of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                               
// AXI_EXOKAY_RESPONSE_NORMAL_READ                                             -  60072 -  Slave has responded ~AXI_EXOKAY~ to a non exclusive read transfer                                                                                                                
// AXI_EXOKAY_RESPONSE_NORMAL_WRITE                                            -  60073 -  Slave has responded ~AXI_EXOKAY~ to a non exclusive write transfer                                                                                                               
// AXI_EX_RD_RESP_MISMATCHED_WITH_EXPECTED_RESP                                -  60074 -  Expected response to this exclusive read did not matched with the actual response (SPEC3(A7.2.3))                                                                            
// AXI_EX_WR_RESP_MISMATCHED_WITH_EXPECTED_RESP                                -  60075 -  Expected response to this exclusive write did not matched with the actual response (SPEC3(A7.2.3))                                                                           
// AXI_EX_RD_EXOKAY_RESP_SLAVE_WITHOUT_EXCLUSIVE_ACCESS                        -  60076 -  Response for an exclusive read to a slave which does not support exclusive access should be ~AXI_OKAY~, but it returned ~AXI_EXOKAY~ (SPEC3(A7.2.3))
// AXI_EX_WRITE_BEFORE_EX_READ_RESPONSE                                        -  60077 -  Exclusive write has occurred, with no previous exclusive read (SPEC3(A7.2.2))                                                                                                        
// AXI_EX_WRITE_EXOKAY_RESP_SLAVE_WITHOUT_EXCLUSIVE_ACCESS                     -  60078 -  Response for an exclusive write to a slave which does not support exclusive access should be ~AXI_OKAY~, but it returned ~AXI_EXOKAY~ (SPEC3(A7.2.3))              
// AXI_ILLEGAL_LENGTH_WRAPPING_READ_BURST                                      -  60079 -  In the last read address phase burst_length has an illegal value for a burst of type AXI_WRAP (SPEC3(A3.4.1))                                                         
// AXI_ILLEGAL_LENGTH_WRAPPING_WRITE_BURST                                     -  60080 -  In the last write address phase burst_length has an illegal value for a burst of type AXI_WRAP (SPEC3(A3.4.1))                                                        
// AXI_ILLEGAL_RESPONSE_EXCLUSIVE_READ                                         -  60081 -  Response for an exclusive read should be either ~AXI_OKAY~ or ~AXI_EXOKAY~ (SPEC3(A7.2.3))                                                                                    
// AXI_ILLEGAL_RESPONSE_EXCLUSIVE_WRITE                                        -  60082 -  Response for an exclusive write should be either ~AXI_OKAY~ or ~AXI_EXOKAY~ (SPEC3(A7.2.3))                                                                                   
// AXI_PARAM_READ_DATA_BUS_WIDTH                                               -  60083 -  The value of <AXI_RDATA_WIDTH> must be one of 8,16,32,64,128,256,512,1024 (SPEC3(A1.3.1))                                                                                            
// AXI_PARAM_WRITE_DATA_BUS_WIDTH                                              -  60084 -  The value of <AXI_WDATA_WIDTH> must be one of 8,16,32,64,128,256,512,1024 (SPEC3(A1.3.1))                                                                                        
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_12                                    -  60085 -  The RA bit of the cache parameter should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                              
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_13                                    -  60086 -  The RA bit of the cache parameter should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                             
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_4                                     -  60087 -  The RA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                                
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_5                                     -  60088 -  The RA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                                  
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_8                                     -  60089 -  The RA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                                     
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_9                                     -  60090 -  The RA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                                     
// AXI_READ_BURST_LENGTH_VIOLATION                                             -  60091 -  The burst_length implied by the number of beats actually read does not match the burst_length defined by the <axi_master_read_addr_channel_phase> (SPEC3(A3.4.1))                             
// AXI_READ_BURST_SIZE_VIOLATION                                               -  60092 -  In this read transaction, size has been set greater than the defined data bus width (SPEC3(A3.4.1))                                                                                                   
// AXI_READ_DATA_BEFORE_ADDRESS                                                -  60093 -  An unexpected read response has occurred (there are no outstanding read transactions with this id) (SPEC3(A3.3.1))                                                                           
// AXI_READ_DATA_CHANGED_BEFORE_RREADY                                         -  60094 -  The value of <RDATA> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                              
// AXI_READ_DATA_UNKN                                                          -  60095 -  <RDATA> has an X value/<RDATA> has a Z value (SPEC3(A2.6))                                                                                                                                     
// AXI_RESERVED_ARLOCK_ENCODING                                                -  60096 -  The reserved encoding of 2'b11 should not be used for ARLOCK (SPEC3(A7.4))                                                                                                                   
// AXI_READ_RESP_CHANGED_BEFORE_RREADY                                         -  60097 -  The value of <RRESP> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                        
// AXI_RESERVED_ARBURST_ENCODING                                               -  60098 -  The reserved encoding of 2'b11 should not be used for <ARBURST> (SPEC3(A3.4.1))                                                                                              
// AXI_RESERVED_AWBURST_ENCODING                                               -  60099 -  The reserved encoding of 2'b11 should not be used for <AWBURST> (SPEC3(A3.4.1))                                                                                                  
// AXI_RID_CHANGED_BEFORE_RREADY                                               -  60100 -  The value of <RID> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                              
// AXI_RID_UNKN                                                                -  60101 -  <RID> has an X value/<RID> has a Z value (SPEC3(A2.6))                                                                                                                                    
// AXI_RLAST_CHANGED_BEFORE_RREADY                                             -  60102 -  The value of <RLAST> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                     
// AXI_RLAST_UNKN                                                              -  60103 -  <RLAST> has an X value/<RLAST> has a Z value (SPEC3(A2.6))                                                                                                                                 
// AXI_RREADY_UNKN                                                             -  60104 -  <RREADY> has an X value/<RREADY> has a Z value (SPEC3(A2.6))                                                                                                                                   
// AXI_RRESP_UNKN                                                              -  60105 -  <RRESP> has an X value/<RRESP> has a Z value (SPEC3(A2.6))                                                                                                                                  
// AXI_RUSER_CHANGED_BEFORE_RREADY                                             -  60106 -  The value of <RUSER> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                          
// AXI_RUSER_UNKN                                                              -  60107 -  <RUSER> has an X value/<RUSER> has a Z value (SPEC3(A2.6))                                                                                                              
// AXI_RVALID_DEASSERTED_BEFORE_RREADY                                         -  60108 -  <RVALID> has been de-asserted before <RREADY> was asserted (SPEC3(A3.2.1))                                                                         
// AXI_RVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  -  60109 -  A slave interface must begin driving  <RVALID> high only at a rising clock edge after ARESETn is HIGH (SPEC3(A3.1.2))                                  
// AXI_RVALID_UNKN                                                             -  60110 -  <RVALID> has an X value/<RVALID> has a Z value (SPEC3(A2.6))                                                                                                        
// AXI_UNALIGNED_ADDRESS_FOR_EXCLUSIVE_READ                                    -  60111 -  Exclusive read accesses must have address aligned to the total number of bytes in the transaction (SPEC3(A7.2.4))                                     
// AXI_UNALIGNED_ADDRESS_FOR_EXCLUSIVE_WRITE                                   -  60112 -  Exclusive write accesses must have address aligned to the total number of bytes in the transaction (SPEC3(A7.2.4))                                     
// AXI_UNALIGNED_ADDR_FOR_WRAPPING_READ_BURST                                  -  60113 -  Wrapping bursts must have address aligned to the start of the read transfer (SPEC3(A3.4.1))                                                                                                                                    
// AXI_UNALIGNED_ADDR_FOR_WRAPPING_WRITE_BURST                                 -  60114 -  Wrapping bursts must have address aligned to the start of the write transfet (SPEC3(A3.4.1))                                                                                                                                    
// AXI_WDATA_CHANGED_BEFORE_WREADY_ON_INVALID_LANE                             -  60115 -  On a lane whose strobe is 0, the value of <WDATA> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                               
// AXI_WDATA_CHANGED_BEFORE_WREADY_ON_VALID_LANE                               -  60116 -  On a lane whose strobe is 1, the value of <WDATA> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                   
// AXI_WLAST_CHANGED_BEFORE_WREADY                                             -  60117 -  The value of <WLAST> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                
// AXI_WID_CHANGED_BEFORE_WREADY                                               -  60118 -  The value of <WID> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                
// AXI_WLAST_UNKN                                                              -  60119 -  <WLAST> has an X value/<WLAST> has an Z value (SPEC3(A2.3))                                                                                        
// AXI_WID_UNKN                                                                -  60120 -  <WID> has an X value/<WID> has an Z value (SPEC3(A2.3))                                                                                                     
// AXI_WREADY_UNKN                                                             -  60121 -  <WREADY> has an X value/<WREADY> has a Z value (SPEC3(A2.3))                                                                                       
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_12                                   -  60122 -  The WA bit of the cache parameter should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                     
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_13                                   -  60123 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                   
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_4                                    -  60124 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                              
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_5                                    -  60125 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                         
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_8                                    -  60126 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                           
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_9                                    -  60127 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                            
// AXI_WRITE_BURST_SIZE_VIOLATION                                              -  60128 -  In this write transaction, size has been set greater than the defined data buswidth (SPEC3(A3.4.1))                                         
// AXI_WRITE_DATA_BEFORE_ADDRESS                                               -  60129 -  A write data beat has occurred before the corresponding address phase                                                                      
// AXI_WRITE_DATA_UNKN_ON_INVALID_LANE                                         -  60130 -  DEPRECATED - This assertion is now DEPRECATED and by default DISABLED, as per protocol Byte lanes for which strobe is 0 could take unknown value..
// AXI_WRITE_DATA_UNKN_ON_VALID_LANE                                           -  60131 -  On a lane whose strobe is 1, <WDATA> has an X value/<WDATA> has a Z value (SPEC3(A2.3))                                          
// AXI_RESERVED_AWLOCK_ENCODING                                                -  60132 -  The reserved encoding of 2'b11 should not be used for AWLOCK (SPEC3(A7.4))                                                                                                                                
// AXI_WRITE_STROBE_ON_INVALID_BYTE_LANES                                      -  60133 -  Write strobe(s) incorrect for the address/size of a fixed transfer (SPEC3(A2.3))                                                                                                                  
// AXI_WSTRB_CHANGED_BEFORE_WREADY                                             -  60134 -  The value of <WSTRB> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                         
// AXI_WSTRB_UNKN                                                              -  60135 -  <WSTRB> has an X value/<WSTRB> has an Z value (SPEC3(A2.3))                                                                                                                                                      
// AXI_WUSER_CHANGED_BEFORE_WREADY                                             -  60136 -  The value of <WUSER> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                        
// AXI_WUSER_UNKN                                                              -  60137 -  <WUSER> has an X value/<WUSER> has an Z value (SPEC3(A2.3))                                                                                                                              
// AXI_WVALID_DEASSERTED_BEFORE_WREADY                                         -  60138 -  <WVALID> has been de-asserted before <WREADY> was asserted (SPEC3(A3.2.1))                                                                                               
// AXI_WVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  -  60139 -  A master interface must begin driving <WVALID> high only at a rising clock edge after <ARESETn> is HIGH (SPEC3(A3.1.2))                                             
// AXI_WVALID_UNKN                                                             -  60140 -  <WVALID> has an X value/<WVALID> has an Z value (SPEC3(A2.3))                                                                                                             
// AXI_ADDR_ACROSS_4K_WITHIN_LOCKED_WRITE_TRANSACTION                          -  60141 -  Transactions within a locked write sequence should be within the same 4K address boundary (SPEC3(A7.3))                                           
// AXI_ADDR_ACROSS_4K_WITHIN_LOCKED_READ_TRANSACTION                           -  60142 -  Transactions within a locked read sequence should be within the same 4K address boundary (SPEC3(A7.3))                                            
// AXI_AWID_CHANGED_WITHIN_LOCKED_TRANSACTION                                  -  60143 -  Master should not change the awid within the locked transaction (SPEC3(A7.3))                                               
// AXI_ARID_CHANGED_WITHIN_LOCKED_TRANSACTION                                  -  60144 -  Master should not change the arid within the locked transaction (SPEC3(A7.3))                                              
// AXI_AWPROT_CHANGED_WITHIN_LOCKED_TRANSACTION                                -  60145 -  Master should not change the awprot within the locked transaction (SPEC3(A7.3))                                                   
// AXI_ARPROT_CHANGED_WITHIN_LOCKED_TRANSACTION                                -  60146 -  Master should not change the arprot within the locked transaction (SPEC3(A7.3))                                                 
// AXI_AWCACHE_CHANGED_WITHIN_LOCKED_TRANSACTION                               -  60147 -  Master should not change the awcache within the locked transaction (SPEC3(A7.3))                                                    
// AXI_ARCACHE_CHANGED_WITHIN_LOCKED_TRANSACTION                               -  60148 -  Master should not change the arcache within the locked transaction (SPEC3(A7.3))                                                      
// AXI_NUMBER_OF_LOCKED_SEQUENCES_EXCEEDS_2                                    -  60149 -  Number of accesses within a locked sequence should not be more than 2 (SPEC3(A7.3))                                                                                                     
// AXI_LOCKED_WRITE_BEFORE_COMPLETION_OF_PREVIOUS_WRITE_TRANSACTIONS           -  60150 -  A locked write sequence should not commence before completion of all previously issued write addresses (SPEC3(A7.3))                                                 
// AXI_LOCKED_WRITE_BEFORE_COMPLETION_OF_PREVIOUS_READ_TRANSACTIONS            -  60151 -  A locked write sequence should not commence before completion of all previously issued read addresses (SPEC3(A7.3))                                              
// AXI_LOCKED_READ_BEFORE_COMPLETION_OF_PREVIOUS_WRITE_TRANSACTIONS            -  60152 -  A locked read sequence should not commence before completion of all previously issued write addresses (SPEC3(A7.3))                                                    
// AXI_LOCKED_READ_BEFORE_COMPLETION_OF_PREVIOUS_READ_TRANSACTIONS             -  60153 -  A locked read sequence should not commence before completion of all previously issued read addresses (SPEC3(A7.3))                                                        
// AXI_NEW_BURST_BEFORE_COMPLETION_OF_UNLOCK_TRANSACTION                       -  60154 -  The unlocking transaction should be completed before further any transactions are initiated (SPEC3(A7.3))                                                           
// AXI_UNLOCKED_WRITE_WHILE_OUTSTANDING_LOCKED_WRITES                          -  60155 -  Unlocking write transaction started while outstanding locked write transaction has not completed (SPEC3(A7.3))                                                  
// AXI_UNLOCKED_WRITE_WHILE_OUTSTANDING_LOCKED_READS                           -  60156 -  Unlocking write transaction started while outstanding locked read transaction has not completed (SPEC3(A7.3))                                                 
// AXI_UNLOCKED_READ_WHILE_OUTSTANDING_LOCKED_WRITES                           -  60157 -  Unlocking read transaction started while outstanding locked write transaction has not completed (SPEC3(A7.3))                                                             
// AXI_UNLOCKED_READ_WHILE_OUTSTANDING_LOCKED_READS                            -  60158 -  Unlocking read transaction started while outstanding locked read transaction has not completed (SPEC3(A7.3))                                                     
// AXI_UNLOCKING_TRANSACTION_WITH_AN_EXCLUSIVE_ACCESS                          -  60159 -  Unlocking transaction can not be an exclusive access transaction (SPEC3(A7.3))                                                                                                                                                            
// AXI_FIRST_DATA_ITEM_OF_TRANSACTION_WRITE_ORDER_VIOLATION                    -  60160 -  The order in which a slave receives the first data item of each transaction must be the same as the order in which it receives the addresses for the transaction (SPEC3(A5.3.3))                                                      
// AXI_AWLEN_MISMATCHED_WITH_COMPLETED_WRITE_DATA_BURST                        -  60161 -  AWLEN value of write address control does not match with corresponding outstanding write data burts length (SPEC3(A3.4.1))                                                       
// AXI_WRITE_LENGTH_MISMATCHED_ACTUAL_LENGTH_OF_WRITE_DATA_BURST_EXCEEDS_AWLEN -  60162 -  The actual length of write data burst exceeds with the length specified by AWLEN (SPEC3(A3.4.1))                                              
// AXI_AWLEN_MISMATCHED_ACTUAL_LENGTH_OF_WRITE_DATA_BURST_EXCEEDS_AWLEN        -  60163 -  Actual length of data burst has exceeded the burst length specified by AWLEN (SPEC3(A3.4.1))                                                               
// AXI_WLAST_ASSERTED_DURING_DATA_PHASE_OTHER_THAN_LAST                        -  60164 -  AWLEN value of write address control does not match with corresponding outstanding write data burts length (SPEC3(A3.4.1))                                                 
// AXI_WRITE_INTERLEAVE_DEPTH_VIOLATION                                        -  60165 -  Write data bursts should not be interleaved beyond the write interleaving depth (SPEC3(A5.3.3))                                   
// AXI_WRITE_RESPONSE_WITHOUT_ADDR                                             -  60166 -  Write response should not be sent before the corresponding address has completed (SPEC3(A3.3.1))                                 
// AXI_WRITE_RESPONSE_WITHOUT_DATA                                             -  60167 -  Write response should not be sent before the corresponding write data burst completed (SPEC3(A3.3.1))                           
// AXI_AWVALID_HIGH_DURING_RESET                                               -  60168 -  AWVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                     
// AXI_WVALID_HIGH_DURING_RESET                                                -  60169 -  WVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                       
// AXI_BVALID_HIGH_DURING_RESET                                                -  60170 -  BVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                        
// AXI_ARVALID_HIGH_DURING_RESET                                               -  60171 -  ARVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                          
// AXI_RVALID_HIGH_DURING_RESET                                                -  60172 -  RVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                         
// AXI_RLAST_VIOLATION                                                         -  60173 -  RLAST signal should be asserted along with the final transfer of the read data burst (SPEC3(A3.4.1))                                                                                    
// AXI_EX_WRITE_AFTER_EX_READ_FAILURE                                          -  60174 -  It is recommended that an exclusive write access should not be performed after the corresponding exclusive read failure. (SPEC3(A7.2.2))                                
// AXI_TIMEOUT_WAITING_FOR_WRITE_DATA                                          -  60175 -  Timed-out waiting for a data phase in write data burst. SPEC3(A2.3)                                                           
// AXI_TIMEOUT_WAITING_FOR_WRITE_RESPONSE                                      -  60176 -  Timed-out waiting for a write response. SPEC3(A2.4)                                                                      
// AXI_TIMEOUT_WAITING_FOR_READ_RESPONSE                                       -  60177 -  Timed-out waiting for a read response. SPEC3(A2.6)                                                                            
// AXI_TIMEOUT_WAITING_FOR_WRITE_ADDR_AFTER_DATA                               -  60178 -  Timed-out waiting for a write address phase to be coming after data SPEC3(A2.2)                                       
// AXI_DEC_ERR_RESP_FOR_READ                                                   -  60179 -  No slave at the address for this read transfer (signaled by ~AXI_DECERR~)                                                                     
// AXI_DEC_ERR_RESP_FOR_WRITE                                                  -  60180 -  No slave at the address for this write transfer (signaled by ~AXI_DECERR~)                                                                     
// AXI_SLV_ERR_RESP_FOR_READ                                                   -  60181 -  Slave has detected an error for this read transfer (signaled by ~AXI_SLVERR~)                                                                  
// AXI_SLV_ERR_RESP_FOR_WRITE                                                  -  60182 -  Slave has detected an error for this write transfer (signaled by ~AXI_SLVERR~)                                                                   
// AXI_MINIMUM_SLAVE_ADDRESS_SPACE_VIOLATION                                   -  60183 -  The minimum address space occupied by a single slave device is 4 kilobytes (SPEC3(A10.3.2))                                       
// AXI_ADDRESS_WIDTH_EXCEEDS_64                                                -  60184 -  AXI supports up to 64-bit addressing (SPEC3(A10.3.1))                                                                                                                  
// AXI_READ_BURST_MAXIMUM_LENGTH_VIOLATION                                     -  60185 -  16 read data beats were seen without RLAST (SPEC3(A3.4.1))                                                                                                   
// AXI_WRITE_BURST_MAXIMUM_LENGTH_VIOLATION                                    -  60186 -  16 write data beats were seen without WLAST (see AMBA AXI and ACE Protocol Specification IHI0022D section A3.4.1 )                                     
// AXI_WRITE_STROBES_LENGTH_VIOLATION                                          -  60187 -  The size of the write_strobes array in a write transfer should match the value given by AWLEN                                                                                               
// AXI_EX_RD_WHEN_EX_NOT_ENABLED                                               -  60188 -  An exclusive read should not be issued when exclusive transactions are not enabled                                                                                                                   
// AXI_EX_WR_WHEN_EX_NOT_ENABLED                                               -  60189 -  An exclusive write should not be issued when exclusive transactions are not enabled                                                                                                     
// AXI_WRITE_TRANSFER_EXCEEDS_ADDRESS_SPACE                                    -  60190 -  This write transfer runs off the edge of the address space defined by AXI_ADDRESS_WIDTH (SPEC3(A10.3.1))                                                                           
// AXI_READ_TRANSFER_EXCEEDS_ADDRESS_SPACE                                     -  60191 -  This read transfer runs off the edge of the address space defined by AXI_ADDRESS_WIDTH (SPEC3(A10.3.1))                                                                                 
// AXI_EXCL_RD_WHILE_EXCL_WR_IN_PROGRESS_SAME_ID                               -  60192 -  Master starts an exclusive read burst while exclusive write burst with same ID tag is in progress (SPEC3(A7.2.4))                                                                 
// AXI_EXCL_WR_WHILE_EXCL_RD_IN_PROGRESS_SAME_ID                               -  60193 -  Master starts an exclusive write burst while exclusive read burst with same ID tag is in progress (SPEC3(A7.2.4))                                                                
// AXI_ILLEGAL_LENGTH_READ_BURST                                               -  60194 -  Read address phase burst_length has an illegal value (SPEC3(A3.4.1))                                                                                                                      
// AXI_ILLEGAL_LENGTH_WRITE_BURST                                              -  60195 -  Write address phase burst_length has an illegal value (SPEC3(A3.4.1))                                                                                                                        
// AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID                                      -  60196 -  Once ARVALID has been asserted, ARREADY> should be asserted within config_max_latency_ARVALID_assertion_to_ARREADY clock periods                                                     
// AXI_BREADY_NOT_ASSERTED_AFTER_BVALID                                        -  60197 -  Once BVALID has been asserted, BREADY> should be asserted within config_max_latency_BVALID_assertion_to_BREADY clock periods                                                             
// AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID                                      -  60198 -  Once AWVALID has been asserted, AWREADY> should be asserted within config_max_latency_AWVALID_assertion_to_AWREADY clock periods                                                              
// AXI_RREADY_NOT_ASSERTED_AFTER_RVALID                                        -  60199 -  Once RVALID has been asserted, RREADY> should be asserted within config_max_latency_RVALID_assertion_to_RREADY clock periods                                                                
// AXI_WREADY_NOT_ASSERTED_AFTER_WVALID                                        -  60200 -  Once WVALID has been asserted, WREADY> should be asserted within config_max_latency_WVALID_assertion_to_WREADY clock periods                                                           
// AXI_DEC_ERR_ILLEGAL_FOR_MAPPED_SLAVE_ADDR                                   -  60201 -  Slave receives a burst to a mapped address but responds with DECERR (signalled by AXI_DECERR) (SPEC3(A3.4.4))                                                                           
// AXI_PARAM_READ_REORDERING_DEPTH_EQUALS_ZERO                                 -  60202 -  The user-supplied config_read_data_reordering_depth should be greater than zero (SPEC3(A5.3.1))                                                                                        
// AXI_PARAM_READ_REORDERING_DEPTH_EXCEEDS_MAX_ID                              -  60203 -  The user-supplied config_read_data_reordering_depth exceeds the maximum possible value, as defined by the AXI_ID_WIDTH parameter (SPEC3(A5.3.1))                              
// AXI_READ_REORDERING_VIOLATION                                               -  60204 -  The arrival of a read response has exceeded the read reordering depth (SPEC3(A5.3.1))                             
// AXI_READ_ISSUING_CAPABILITY_VIOLATION                                       -  60205 -  Number of outstanding Read transactions exceeded maximum Read issuing capability 
// AXI_WRITE_ISSUING_CAPABILITY_VIOLATION                                      -  60206 -  Number of outstanding Write transactions exceeded maximum Write issuing capability
// AXI_COMBINED_ISSUING_CAPABILITY_VIOLATION                                   -  60207 -  Number of outstanding Read and Write transactions exceeded maximum combined issuing capability 
// AXI_READ_ACCEPTANCE_CAPABILITY_VIOLATION                                    -  60208 -  Number of outstanding Read transactions exceeded maximum Read acceptance capability 
// AXI_WRITE_ACCEPTANCE_CAPABILITY_VIOLATION                                   -  60209 -  Number of outstanding Write transactions exceeded maximum Write acceptance capability 
// AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION                                -  60210 -  Number of outstanding Read and Write transactions exceeded maximum combined acceptance capability 
typedef enum bit [7:0]
{
    AXI_ARESETn_SIGNAL_Z                                                        = 8'h00,
    AXI_ARESETn_SIGNAL_X                                                        = 8'h01,
    AXI_ACLK_SIGNAL_Z                                                           = 8'h02,
    AXI_ACLK_SIGNAL_X                                                           = 8'h03,
    AXI_ADDR_FOR_READ_BURST_ACROSS_4K_BOUNDARY                                  = 8'h04,
    AXI_ADDR_FOR_WRITE_BURST_ACROSS_4K_BOUNDARY                                 = 8'h05,
    AXI_ARADDR_CHANGED_BEFORE_ARREADY                                           = 8'h06,
    AXI_ARADDR_UNKN                                                             = 8'h07,
    AXI_ARBURST_CHANGED_BEFORE_ARREADY                                          = 8'h08,
    AXI_ARBURST_UNKN                                                            = 8'h09,
    AXI_ARCACHE_CHANGED_BEFORE_ARREADY                                          = 8'h0a,
    AXI_ARCACHE_UNKN                                                            = 8'h0b,
    AXI_ARID_CHANGED_BEFORE_ARREADY                                             = 8'h0c,
    AXI_ARID_UNKN                                                               = 8'h0d,
    AXI_ARLEN_CHANGED_BEFORE_ARREADY                                            = 8'h0e,
    AXI_ARLEN_UNKN                                                              = 8'h0f,
    AXI_ARLOCK_CHANGED_BEFORE_ARREADY                                           = 8'h10,
    AXI_ARLOCK_UNKN                                                             = 8'h11,
    AXI_ARPROT_CHANGED_BEFORE_ARREADY                                           = 8'h12,
    AXI_ARPROT_UNKN                                                             = 8'h13,
    AXI_ARREADY_UNKN                                                            = 8'h14,
    AXI_ARSIZE_CHANGED_BEFORE_ARREADY                                           = 8'h15,
    AXI_ARSIZE_UNKN                                                             = 8'h16,
    AXI_ARUSER_CHANGED_BEFORE_ARREADY                                           = 8'h17,
    AXI_ARUSER_UNKN                                                             = 8'h18,
    AXI_ARVALID_DEASSERTED_BEFORE_ARREADY                                       = 8'h19,
    AXI_ARVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                 = 8'h1a,
    AXI_ARVALID_UNKN                                                            = 8'h1b,
    AXI_AWADDR_CHANGED_BEFORE_AWREADY                                           = 8'h1c,
    AXI_AWADDR_UNKN                                                             = 8'h1d,
    AXI_AWBURST_CHANGED_BEFORE_AWREADY                                          = 8'h1e,
    AXI_AWBURST_UNKN                                                            = 8'h1f,
    AXI_AWCACHE_CHANGED_BEFORE_AWREADY                                          = 8'h20,
    AXI_AWCACHE_UNKN                                                            = 8'h21,
    AXI_AWID_CHANGED_BEFORE_AWREADY                                             = 8'h22,
    AXI_AWID_UNKN                                                               = 8'h23,
    AXI_AWLEN_CHANGED_BEFORE_AWREADY                                            = 8'h24,
    AXI_AWLEN_UNKN                                                              = 8'h25,
    AXI_AWLOCK_CHANGED_BEFORE_AWREADY                                           = 8'h26,
    AXI_AWLOCK_UNKN                                                             = 8'h27,
    AXI_AWPROT_CHANGED_BEFORE_AWREADY                                           = 8'h28,
    AXI_AWPROT_UNKN                                                             = 8'h29,
    AXI_AWREADY_UNKN                                                            = 8'h2a,
    AXI_AWSIZE_CHANGED_BEFORE_AWREADY                                           = 8'h2b,
    AXI_AWSIZE_UNKN                                                             = 8'h2c,
    AXI_AWUSER_CHANGED_BEFORE_AWREADY                                           = 8'h2d,
    AXI_AWUSER_UNKN                                                             = 8'h2e,
    AXI_AWVALID_DEASSERTED_BEFORE_AWREADY                                       = 8'h2f,
    AXI_AWVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                 = 8'h30,
    AXI_AWVALID_UNKN                                                            = 8'h31,
    AXI_BID_CHANGED_BEFORE_BREADY                                               = 8'h32,
    AXI_BID_UNKN                                                                = 8'h33,
    AXI_BREADY_UNKN                                                             = 8'h34,
    AXI_BRESP_CHANGED_BEFORE_BREADY                                             = 8'h35,
    AXI_BRESP_UNKN                                                              = 8'h36,
    AXI_BUSER_CHANGED_BEFORE_BREADY                                             = 8'h37,
    AXI_BUSER_UNKN                                                              = 8'h38,
    AXI_BVALID_DEASSERTED_BEFORE_BREADY                                         = 8'h39,
    AXI_BVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  = 8'h3a,
    AXI_BVALID_UNKN                                                             = 8'h3b,
    AXI_EXCLUSIVE_READ_ACCESS_MODIFIABLE                                        = 8'h3c,
    AXI_EXCLUSIVE_READ_BYTES_TRANSFER_EXCEEDS_128                               = 8'h3d,
    AXI_EXCLUSIVE_WRITE_BYTES_TRANSFER_EXCEEDS_128                              = 8'h3e,
    AXI_EXCLUSIVE_READ_BYTES_TRANSFER_NOT_POWER_OF_2                            = 8'h3f,
    AXI_EXCLUSIVE_WRITE_BYTES_TRANSFER_NOT_POWER_OF_2                           = 8'h40,
    AXI_EXCLUSIVE_WR_ADDRESS_NOT_SAME_AS_RD                                     = 8'h41,
    AXI_EXCLUSIVE_WR_BURST_NOT_SAME_AS_RD                                       = 8'h42,
    AXI_EXCLUSIVE_WR_CACHE_NOT_SAME_AS_RD                                       = 8'h43,
    AXI_EXCLUSIVE_WRITE_ACCESS_MODIFIABLE                                       = 8'h44,
    AXI_EXCLUSIVE_WR_LENGTH_NOT_SAME_AS_RD                                      = 8'h45,
    AXI_EXCLUSIVE_WR_PROT_NOT_SAME_AS_RD                                        = 8'h46,
    AXI_EXCLUSIVE_WR_SIZE_NOT_SAME_AS_RD                                        = 8'h47,
    AXI_EXOKAY_RESPONSE_NORMAL_READ                                             = 8'h48,
    AXI_EXOKAY_RESPONSE_NORMAL_WRITE                                            = 8'h49,
    AXI_EX_RD_RESP_MISMATCHED_WITH_EXPECTED_RESP                                = 8'h4a,
    AXI_EX_WR_RESP_MISMATCHED_WITH_EXPECTED_RESP                                = 8'h4b,
    AXI_EX_RD_EXOKAY_RESP_SLAVE_WITHOUT_EXCLUSIVE_ACCESS                        = 8'h4c,
    AXI_EX_WRITE_BEFORE_EX_READ_RESPONSE                                        = 8'h4d,
    AXI_EX_WRITE_EXOKAY_RESP_SLAVE_WITHOUT_EXCLUSIVE_ACCESS                     = 8'h4e,
    AXI_ILLEGAL_LENGTH_WRAPPING_READ_BURST                                      = 8'h4f,
    AXI_ILLEGAL_LENGTH_WRAPPING_WRITE_BURST                                     = 8'h50,
    AXI_ILLEGAL_RESPONSE_EXCLUSIVE_READ                                         = 8'h51,
    AXI_ILLEGAL_RESPONSE_EXCLUSIVE_WRITE                                        = 8'h52,
    AXI_PARAM_READ_DATA_BUS_WIDTH                                               = 8'h53,
    AXI_PARAM_WRITE_DATA_BUS_WIDTH                                              = 8'h54,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_12                                    = 8'h55,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_13                                    = 8'h56,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_4                                     = 8'h57,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_5                                     = 8'h58,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_8                                     = 8'h59,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_9                                     = 8'h5a,
    AXI_READ_BURST_LENGTH_VIOLATION                                             = 8'h5b,
    AXI_READ_BURST_SIZE_VIOLATION                                               = 8'h5c,
    AXI_READ_DATA_BEFORE_ADDRESS                                                = 8'h5d,
    AXI_READ_DATA_CHANGED_BEFORE_RREADY                                         = 8'h5e,
    AXI_READ_DATA_UNKN                                                          = 8'h5f,
    AXI_RESERVED_ARLOCK_ENCODING                                                = 8'h60,
    AXI_READ_RESP_CHANGED_BEFORE_RREADY                                         = 8'h61,
    AXI_RESERVED_ARBURST_ENCODING                                               = 8'h62,
    AXI_RESERVED_AWBURST_ENCODING                                               = 8'h63,
    AXI_RID_CHANGED_BEFORE_RREADY                                               = 8'h64,
    AXI_RID_UNKN                                                                = 8'h65,
    AXI_RLAST_CHANGED_BEFORE_RREADY                                             = 8'h66,
    AXI_RLAST_UNKN                                                              = 8'h67,
    AXI_RREADY_UNKN                                                             = 8'h68,
    AXI_RRESP_UNKN                                                              = 8'h69,
    AXI_RUSER_CHANGED_BEFORE_RREADY                                             = 8'h6a,
    AXI_RUSER_UNKN                                                              = 8'h6b,
    AXI_RVALID_DEASSERTED_BEFORE_RREADY                                         = 8'h6c,
    AXI_RVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  = 8'h6d,
    AXI_RVALID_UNKN                                                             = 8'h6e,
    AXI_UNALIGNED_ADDRESS_FOR_EXCLUSIVE_READ                                    = 8'h6f,
    AXI_UNALIGNED_ADDRESS_FOR_EXCLUSIVE_WRITE                                   = 8'h70,
    AXI_UNALIGNED_ADDR_FOR_WRAPPING_READ_BURST                                  = 8'h71,
    AXI_UNALIGNED_ADDR_FOR_WRAPPING_WRITE_BURST                                 = 8'h72,
    AXI_WDATA_CHANGED_BEFORE_WREADY_ON_INVALID_LANE                             = 8'h73,
    AXI_WDATA_CHANGED_BEFORE_WREADY_ON_VALID_LANE                               = 8'h74,
    AXI_WLAST_CHANGED_BEFORE_WREADY                                             = 8'h75,
    AXI_WID_CHANGED_BEFORE_WREADY                                               = 8'h76,
    AXI_WLAST_UNKN                                                              = 8'h77,
    AXI_WID_UNKN                                                                = 8'h78,
    AXI_WREADY_UNKN                                                             = 8'h79,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_12                                   = 8'h7a,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_13                                   = 8'h7b,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_4                                    = 8'h7c,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_5                                    = 8'h7d,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_8                                    = 8'h7e,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_9                                    = 8'h7f,
    AXI_WRITE_BURST_SIZE_VIOLATION                                              = 8'h80,
    AXI_WRITE_DATA_BEFORE_ADDRESS                                               = 8'h81,
    AXI_WRITE_DATA_UNKN_ON_INVALID_LANE                                         = 8'h82,
    AXI_WRITE_DATA_UNKN_ON_VALID_LANE                                           = 8'h83,
    AXI_RESERVED_AWLOCK_ENCODING                                                = 8'h84,
    AXI_WRITE_STROBE_ON_INVALID_BYTE_LANES                                      = 8'h85,
    AXI_WSTRB_CHANGED_BEFORE_WREADY                                             = 8'h86,
    AXI_WSTRB_UNKN                                                              = 8'h87,
    AXI_WUSER_CHANGED_BEFORE_WREADY                                             = 8'h88,
    AXI_WUSER_UNKN                                                              = 8'h89,
    AXI_WVALID_DEASSERTED_BEFORE_WREADY                                         = 8'h8a,
    AXI_WVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  = 8'h8b,
    AXI_WVALID_UNKN                                                             = 8'h8c,
    AXI_ADDR_ACROSS_4K_WITHIN_LOCKED_WRITE_TRANSACTION                          = 8'h8d,
    AXI_ADDR_ACROSS_4K_WITHIN_LOCKED_READ_TRANSACTION                           = 8'h8e,
    AXI_AWID_CHANGED_WITHIN_LOCKED_TRANSACTION                                  = 8'h8f,
    AXI_ARID_CHANGED_WITHIN_LOCKED_TRANSACTION                                  = 8'h90,
    AXI_AWPROT_CHANGED_WITHIN_LOCKED_TRANSACTION                                = 8'h91,
    AXI_ARPROT_CHANGED_WITHIN_LOCKED_TRANSACTION                                = 8'h92,
    AXI_AWCACHE_CHANGED_WITHIN_LOCKED_TRANSACTION                               = 8'h93,
    AXI_ARCACHE_CHANGED_WITHIN_LOCKED_TRANSACTION                               = 8'h94,
    AXI_NUMBER_OF_LOCKED_SEQUENCES_EXCEEDS_2                                    = 8'h95,
    AXI_LOCKED_WRITE_BEFORE_COMPLETION_OF_PREVIOUS_WRITE_TRANSACTIONS           = 8'h96,
    AXI_LOCKED_WRITE_BEFORE_COMPLETION_OF_PREVIOUS_READ_TRANSACTIONS            = 8'h97,
    AXI_LOCKED_READ_BEFORE_COMPLETION_OF_PREVIOUS_WRITE_TRANSACTIONS            = 8'h98,
    AXI_LOCKED_READ_BEFORE_COMPLETION_OF_PREVIOUS_READ_TRANSACTIONS             = 8'h99,
    AXI_NEW_BURST_BEFORE_COMPLETION_OF_UNLOCK_TRANSACTION                       = 8'h9a,
    AXI_UNLOCKED_WRITE_WHILE_OUTSTANDING_LOCKED_WRITES                          = 8'h9b,
    AXI_UNLOCKED_WRITE_WHILE_OUTSTANDING_LOCKED_READS                           = 8'h9c,
    AXI_UNLOCKED_READ_WHILE_OUTSTANDING_LOCKED_WRITES                           = 8'h9d,
    AXI_UNLOCKED_READ_WHILE_OUTSTANDING_LOCKED_READS                            = 8'h9e,
    AXI_UNLOCKING_TRANSACTION_WITH_AN_EXCLUSIVE_ACCESS                          = 8'h9f,
    AXI_FIRST_DATA_ITEM_OF_TRANSACTION_WRITE_ORDER_VIOLATION                    = 8'ha0,
    AXI_AWLEN_MISMATCHED_WITH_COMPLETED_WRITE_DATA_BURST                        = 8'ha1,
    AXI_WRITE_LENGTH_MISMATCHED_ACTUAL_LENGTH_OF_WRITE_DATA_BURST_EXCEEDS_AWLEN = 8'ha2,
    AXI_AWLEN_MISMATCHED_ACTUAL_LENGTH_OF_WRITE_DATA_BURST_EXCEEDS_AWLEN        = 8'ha3,
    AXI_WLAST_ASSERTED_DURING_DATA_PHASE_OTHER_THAN_LAST                        = 8'ha4,
    AXI_WRITE_INTERLEAVE_DEPTH_VIOLATION                                        = 8'ha5,
    AXI_WRITE_RESPONSE_WITHOUT_ADDR                                             = 8'ha6,
    AXI_WRITE_RESPONSE_WITHOUT_DATA                                             = 8'ha7,
    AXI_AWVALID_HIGH_DURING_RESET                                               = 8'ha8,
    AXI_WVALID_HIGH_DURING_RESET                                                = 8'ha9,
    AXI_BVALID_HIGH_DURING_RESET                                                = 8'haa,
    AXI_ARVALID_HIGH_DURING_RESET                                               = 8'hab,
    AXI_RVALID_HIGH_DURING_RESET                                                = 8'hac,
    AXI_RLAST_VIOLATION                                                         = 8'had,
    AXI_EX_WRITE_AFTER_EX_READ_FAILURE                                          = 8'hae,
    AXI_TIMEOUT_WAITING_FOR_WRITE_DATA                                          = 8'haf,
    AXI_TIMEOUT_WAITING_FOR_WRITE_RESPONSE                                      = 8'hb0,
    AXI_TIMEOUT_WAITING_FOR_READ_RESPONSE                                       = 8'hb1,
    AXI_TIMEOUT_WAITING_FOR_WRITE_ADDR_AFTER_DATA                               = 8'hb2,
    AXI_DEC_ERR_RESP_FOR_READ                                                   = 8'hb3,
    AXI_DEC_ERR_RESP_FOR_WRITE                                                  = 8'hb4,
    AXI_SLV_ERR_RESP_FOR_READ                                                   = 8'hb5,
    AXI_SLV_ERR_RESP_FOR_WRITE                                                  = 8'hb6,
    AXI_MINIMUM_SLAVE_ADDRESS_SPACE_VIOLATION                                   = 8'hb7,
    AXI_ADDRESS_WIDTH_EXCEEDS_64                                                = 8'hb8,
    AXI_READ_BURST_MAXIMUM_LENGTH_VIOLATION                                     = 8'hb9,
    AXI_WRITE_BURST_MAXIMUM_LENGTH_VIOLATION                                    = 8'hba,
    AXI_WRITE_STROBES_LENGTH_VIOLATION                                          = 8'hbb,
    AXI_EX_RD_WHEN_EX_NOT_ENABLED                                               = 8'hbc,
    AXI_EX_WR_WHEN_EX_NOT_ENABLED                                               = 8'hbd,
    AXI_WRITE_TRANSFER_EXCEEDS_ADDRESS_SPACE                                    = 8'hbe,
    AXI_READ_TRANSFER_EXCEEDS_ADDRESS_SPACE                                     = 8'hbf,
    AXI_EXCL_RD_WHILE_EXCL_WR_IN_PROGRESS_SAME_ID                               = 8'hc0,
    AXI_EXCL_WR_WHILE_EXCL_RD_IN_PROGRESS_SAME_ID                               = 8'hc1,
    AXI_ILLEGAL_LENGTH_READ_BURST                                               = 8'hc2,
    AXI_ILLEGAL_LENGTH_WRITE_BURST                                              = 8'hc3,
    AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID                                      = 8'hc4,
    AXI_BREADY_NOT_ASSERTED_AFTER_BVALID                                        = 8'hc5,
    AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID                                      = 8'hc6,
    AXI_RREADY_NOT_ASSERTED_AFTER_RVALID                                        = 8'hc7,
    AXI_WREADY_NOT_ASSERTED_AFTER_WVALID                                        = 8'hc8,
    AXI_DEC_ERR_ILLEGAL_FOR_MAPPED_SLAVE_ADDR                                   = 8'hc9,
    AXI_PARAM_READ_REORDERING_DEPTH_EQUALS_ZERO                                 = 8'hca,
    AXI_PARAM_READ_REORDERING_DEPTH_EXCEEDS_MAX_ID                              = 8'hcb,
    AXI_READ_REORDERING_VIOLATION                                               = 8'hcc,
    AXI_READ_ISSUING_CAPABILITY_VIOLATION                                       = 8'hcd,
    AXI_WRITE_ISSUING_CAPABILITY_VIOLATION                                      = 8'hce,
    AXI_COMBINED_ISSUING_CAPABILITY_VIOLATION                                   = 8'hcf,
    AXI_READ_ACCEPTANCE_CAPABILITY_VIOLATION                                    = 8'hd0,
    AXI_WRITE_ACCEPTANCE_CAPABILITY_VIOLATION                                   = 8'hd1,
    AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION                                = 8'hd2
} axi_assertion_e;



//------------------------------------------------------------------------------
//
// Enum: axi_ready_e
//
//------------------------------------------------------------------------------
// 
//  Specifies wait if AXI_NOT_READY and specifies no wait if AXI_READY.
// 
typedef enum bit [0:0]
{
    AXI_NOT_READY = 1'h0,
    AXI_READY     = 1'h1
} axi_ready_e;



//------------------------------------------------------------------------------
//
// Enum: axi_wtrans_phase_e
//
//------------------------------------------------------------------------------
// 
//  An enumerated type used in the coverage collector class
//  <axi_functional_coverage> for encoding the address/data/response type for each
//  phase of a write transaction.
// 
//  As each phase of a write occurs, a field of the <axi_write_trans_record>
//  record is updated with the type (address/data/response) of the phase (this
//  information is used at the end of the transaction to classify the
//  <axi_functional_coverage::axi_wtrans_phase_order_e> phase-ordering type of the
//  transaction).
//  See the <axi_functional_coverage::put_wphase> task.
// 
//  A (ADDR) - The address phase of a write transaction.
//  D (DATA) - The data phase of a write transaction.
//  R (RESP) - The response phase of a write transaction.
// 
typedef enum bit [1:0]
{
    A = 2'h0,
    D = 2'h1,
    R = 2'h2
} axi_wtrans_phase_e;


//------------------------------------------------------------------------------
//
// Struct: axi_rw_txn_counts_s
//
//------------------------------------------------------------------------------

typedef struct packed
{
    int unsigned reads_no_resp;
    int unsigned reads_no_resp_for_id;
    int unsigned waddr_no_resp;
    int unsigned waddr_no_resp_for_id;
    int unsigned wdata_no_resp;
    int unsigned wdata_no_resp_for_id;
    int unsigned writes_no_resp;
    int unsigned writes_no_resp_for_id;
} axi_rw_txn_counts_s;



typedef bit [1023:0] axi_max_bits_t;

// enum: axi_config_e
//
// An enum which fields corresponding to each configuration parameter of the VIP
//    AXI_CONFIG_WRITE_CTRL_TO_DATA_MINTIME - 
//         
//         Sets the delay from start of address phase to start of data phase in a write 
//         transaction (in terms of ACLK).
//         
//         Default: 1 
//         
//         This configuration variable has been deprecated and is maintained 
//         for backward compatibility. However, you can use ~write_address_to_data_delay~ 
//         configuration variable to control the delay between a write address phase 
//         and a write data phase.
//         
//    AXI_CONFIG_ENABLE_ALL_ASSERTIONS - 
//         
//         Enables all protocol assertions. 
//         
//         Default: 1
//         
//    AXI_CONFIG_ENABLE_ASSERTION - 
//         
//         Enables individual protocol assertion.
//         This variable controls whether specific assertion within QVIP (of type <axi_assertion_e>) is enabled or disabled.
//         Individual assertion can be disabled as follows:-
//         //-----------------------------------------------------------------------
//         // < BFM interface>.set_config_enable_assertion_index1(<name of assertion>,1'b0);
//         //-----------------------------------------------------------------------
//         
//         For example, the assertion AXI_READ_DATA_UNKN is disabled as follows:
//         <bfm>.set_config_enable_assertion_index1(AXI_READ_DATA_UNKN, 1'b0); 
//         
//         Here bfm is the AXI interface instance name for which the assertion to be disabled. 
//         
//         Default: All assertions are enabled
//           
//         
//    AXI_CONFIG_SUPPORT_EXCLUSIVE_ACCESS - 
//         
//         Enables exclusive transactions support for slave.
//         If disabled, every exclusive read/write returns an OKAY response,
//         and exclusive write updates memory. 
//         
//         Default: 1  
//         
//    AXI_CONFIG_READ_DATA_REORDERING_DEPTH - 
//         
//         Sets the maximum number of different read transaction addresses for which read 
//         data(response) can be sent in any order from slave. 
//         
//         Default: 2 ** AXI_ID_WIDTH
//         
//    AXI_CONFIG_MAX_TRANSACTION_TIME_FACTOR - 
//          
//         Sets maximum timeout period (in terms of ACLK) for any complete read or write transaction, which
//         includes time period for all individual phases of transaction. 
//         
//         Default: 100000 clock cycles
//         
//    AXI_CONFIG_TIMEOUT_MAX_DATA_TRANSFER - 
//          
//         Sets maximum number of write data beats in a write data burst. 
//         
//         Default: 1024  
//         
//    AXI_CONFIG_BURST_TIMEOUT_FACTOR - 
//          
//         Sets maximum timeout period (in terms of ACLK) between individual phases of a transaction. 
//         
//         Default: 10000 clock cycles 
//         
//    AXI_CONFIG_MAX_LATENCY_AWVALID_ASSERTION_TO_AWREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of AWVALID to assertion of AWREADY.
//         An error message AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID is generated if AWREADY is not asserted
//         after assertion of AWVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MAX_LATENCY_ARVALID_ASSERTION_TO_ARREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of ARVALID to assertion of ARREADY.
//         An error message AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID is generated if ARREADY is not asserted
//         after assertion of ARVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MAX_LATENCY_RVALID_ASSERTION_TO_RREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of RVALID to assertion of RREADY.
//         An error message AXI_RREADY_NOT_ASSERTED_AFTER_RVALID is generated if RREADY is not asserted
//         after assertion of RVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MAX_LATENCY_BVALID_ASSERTION_TO_BREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of BVALID to assertion of BREADY.
//         An error message AXI_BREADY_NOT_ASSERTED_AFTER_BVALID is generated if BREADY is not asserted
//         after assertion of BVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MAX_LATENCY_WVALID_ASSERTION_TO_WREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of WVALID to assertion of WREADY.
//         An error message AXI_WREADY_NOT_ASSERTED_AFTER_WVALID is generated if WREADY is not asserted
//         after assertion of WVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MASTER_ERROR_POSITION - 
//         
//         Sets type of master error.
//         
//    AXI_CONFIG_SETUP_TIME - 
//         
//         Sets number of simulation time units from the setup time to the active 
//         clock edge of ACLK. The setup time will always be less than the time period
//         of the clock. 
//         
//         Default: 0
//         
//    AXI_CONFIG_HOLD_TIME - 
//         
//         Sets number of simulation time units from the hold time to the active 
//         clock edge of ACLK. 
//         
//         Default: 0
//         
//    AXI_CONFIG_MAX_OUTSTANDING_WR -  Configures maximum possible outstanding Write transactions
//    AXI_CONFIG_MAX_OUTSTANDING_RD -  Configures maximum possible outstanding Read transactions
//    AXI_CONFIG_MAX_OUTSTANDING_RW -  Configures maximum possible outstanding Combined (Read and Write) transactions
//    AXI_CONFIG_IS_ISSUING -  Enables Master component to use "config_max_outstanding_wr/config_max_outstanding_rd/config_max_outstanding_rw" variables for transaction issuing capability when set to true

typedef enum bit [7:0]
{
    AXI_CONFIG_WRITE_CTRL_TO_DATA_MINTIME    = 8'd0,
    AXI_CONFIG_MASTER_WRITE_DELAY            = 8'd1,
    AXI_CONFIG_ENABLE_ALL_ASSERTIONS         = 8'd2,
    AXI_CONFIG_ENABLE_ASSERTION              = 8'd3,
    AXI_CONFIG_SLAVE_START_ADDR              = 8'd4,
    AXI_CONFIG_SLAVE_END_ADDR                = 8'd5,
    AXI_CONFIG_SUPPORT_EXCLUSIVE_ACCESS      = 8'd6,
    AXI_CONFIG_READ_DATA_REORDERING_DEPTH    = 8'd7,
    AXI_CONFIG_MAX_TRANSACTION_TIME_FACTOR   = 8'd8,
    AXI_CONFIG_TIMEOUT_MAX_DATA_TRANSFER     = 8'd9,
    AXI_CONFIG_BURST_TIMEOUT_FACTOR          = 8'd10,
    AXI_CONFIG_MAX_LATENCY_AWVALID_ASSERTION_TO_AWREADY = 8'd11,
    AXI_CONFIG_MAX_LATENCY_ARVALID_ASSERTION_TO_ARREADY = 8'd12,
    AXI_CONFIG_MAX_LATENCY_RVALID_ASSERTION_TO_RREADY = 8'd13,
    AXI_CONFIG_MAX_LATENCY_BVALID_ASSERTION_TO_BREADY = 8'd14,
    AXI_CONFIG_MAX_LATENCY_WVALID_ASSERTION_TO_WREADY = 8'd15,
    AXI_CONFIG_MASTER_ERROR_POSITION         = 8'd16,
    AXI_CONFIG_SETUP_TIME                    = 8'd17,
    AXI_CONFIG_HOLD_TIME                     = 8'd18,
    AXI_CONFIG_MAX_OUTSTANDING_WR            = 8'd19,
    AXI_CONFIG_MAX_OUTSTANDING_RD            = 8'd20,
    AXI_CONFIG_MAX_OUTSTANDING_RW            = 8'd21,
    AXI_CONFIG_IS_ISSUING                    = 8'd22
} axi_config_e;

// enum: axi_vhd_if_e
//
// For VHDL use only
typedef enum int
{
    AXI_VHD_SET_CONFIG                         = 32'd0,
    AXI_VHD_GET_CONFIG                         = 32'd1,
    AXI_VHD_CREATE_WRITE_TRANSACTION           = 32'd2,
    AXI_VHD_CREATE_READ_TRANSACTION            = 32'd3,
    AXI_VHD_SET_ADDR                           = 32'd4,
    AXI_VHD_GET_ADDR                           = 32'd5,
    AXI_VHD_SET_SIZE                           = 32'd6,
    AXI_VHD_GET_SIZE                           = 32'd7,
    AXI_VHD_SET_BURST                          = 32'd8,
    AXI_VHD_GET_BURST                          = 32'd9,
    AXI_VHD_SET_LOCK                           = 32'd10,
    AXI_VHD_GET_LOCK                           = 32'd11,
    AXI_VHD_SET_CACHE                          = 32'd12,
    AXI_VHD_GET_CACHE                          = 32'd13,
    AXI_VHD_SET_PROT                           = 32'd14,
    AXI_VHD_GET_PROT                           = 32'd15,
    AXI_VHD_SET_ID                             = 32'd16,
    AXI_VHD_GET_ID                             = 32'd17,
    AXI_VHD_SET_BURST_LENGTH                   = 32'd18,
    AXI_VHD_GET_BURST_LENGTH                   = 32'd19,
    AXI_VHD_SET_DATA_WORDS                     = 32'd20,
    AXI_VHD_GET_DATA_WORDS                     = 32'd21,
    AXI_VHD_SET_WRITE_STROBES                  = 32'd22,
    AXI_VHD_GET_WRITE_STROBES                  = 32'd23,
    AXI_VHD_SET_RESP                           = 32'd24,
    AXI_VHD_GET_RESP                           = 32'd25,
    AXI_VHD_SET_ADDR_USER                      = 32'd26,
    AXI_VHD_GET_ADDR_USER                      = 32'd27,
    AXI_VHD_SET_READ_OR_WRITE                  = 32'd28,
    AXI_VHD_GET_READ_OR_WRITE                  = 32'd29,
    AXI_VHD_SET_ADDRESS_VALID_DELAY            = 32'd30,
    AXI_VHD_GET_ADDRESS_VALID_DELAY            = 32'd31,
    AXI_VHD_SET_DATA_VALID_DELAY               = 32'd32,
    AXI_VHD_GET_DATA_VALID_DELAY               = 32'd33,
    AXI_VHD_SET_WRITE_RESPONSE_VALID_DELAY     = 32'd34,
    AXI_VHD_GET_WRITE_RESPONSE_VALID_DELAY     = 32'd35,
    AXI_VHD_SET_ADDRESS_READY_DELAY            = 32'd36,
    AXI_VHD_GET_ADDRESS_READY_DELAY            = 32'd37,
    AXI_VHD_SET_DATA_READY_DELAY               = 32'd38,
    AXI_VHD_GET_DATA_READY_DELAY               = 32'd39,
    AXI_VHD_SET_WRITE_RESPONSE_READY_DELAY     = 32'd40,
    AXI_VHD_GET_WRITE_RESPONSE_READY_DELAY     = 32'd41,
    AXI_VHD_SET_GEN_WRITE_STROBES              = 32'd42,
    AXI_VHD_GET_GEN_WRITE_STROBES              = 32'd43,
    AXI_VHD_SET_OPERATION_MODE                 = 32'd44,
    AXI_VHD_GET_OPERATION_MODE                 = 32'd45,
    AXI_VHD_SET_DELAY_MODE                     = 32'd46,
    AXI_VHD_GET_DELAY_MODE                     = 32'd47,
    AXI_VHD_SET_WRITE_DATA_MODE                = 32'd48,
    AXI_VHD_GET_WRITE_DATA_MODE                = 32'd49,
    AXI_VHD_SET_DATA_BEAT_DONE                 = 32'd50,
    AXI_VHD_GET_DATA_BEAT_DONE                 = 32'd51,
    AXI_VHD_SET_TRANSACTION_DONE               = 32'd52,
    AXI_VHD_GET_TRANSACTION_DONE               = 32'd53,
    AXI_VHD_EXECUTE_TRANSACTION                = 32'd54,
    AXI_VHD_GET_RW_TRANSACTION                 = 32'd55,
    AXI_VHD_EXECUTE_READ_DATA_BURST            = 32'd56,
    AXI_VHD_GET_READ_DATA_BURST                = 32'd57,
    AXI_VHD_EXECUTE_WRITE_DATA_BURST           = 32'd58,
    AXI_VHD_GET_WRITE_DATA_BURST               = 32'd59,
    AXI_VHD_EXECUTE_READ_ADDR_PHASE            = 32'd60,
    AXI_VHD_GET_READ_ADDR_PHASE                = 32'd61,
    AXI_VHD_EXECUTE_READ_DATA_PHASE            = 32'd62,
    AXI_VHD_GET_READ_DATA_PHASE                = 32'd63,
    AXI_VHD_EXECUTE_WRITE_ADDR_PHASE           = 32'd64,
    AXI_VHD_GET_WRITE_ADDR_PHASE               = 32'd65,
    AXI_VHD_EXECUTE_WRITE_DATA_PHASE           = 32'd66,
    AXI_VHD_GET_WRITE_DATA_PHASE               = 32'd67,
    AXI_VHD_EXECUTE_WRITE_RESPONSE_PHASE       = 32'd68,
    AXI_VHD_GET_WRITE_RESPONSE_PHASE           = 32'd69,
    AXI_VHD_CREATE_MONITOR_TRANSACTION         = 32'd70,
    AXI_VHD_CREATE_SLAVE_TRANSACTION           = 32'd71,
    AXI_VHD_PUSH_TRANSACTION_ID                = 32'd72,
    AXI_VHD_POP_TRANSACTION_ID                 = 32'd73,
    AXI_VHD_GET_WRITE_ADDR_DATA                = 32'd74,
    AXI_VHD_GET_READ_ADDR                      = 32'd75,
    AXI_VHD_SET_READ_DATA                      = 32'd76,
    AXI_VHD_PRINT                              = 32'd77,
    AXI_VHD_DESTRUCT_TRANSACTION               = 32'd78,
    AXI_VHD_WAIT_ON                            = 32'd79
} axi_vhd_if_e;


typedef enum bit [7:0]
{
    AXI_CLOCK_POSEDGE = 8'd0,
    AXI_CLOCK_NEGEDGE = 8'd1,
    AXI_CLOCK_ANYEDGE = 8'd2,
    AXI_CLOCK_0_TO_1  = 8'd3,
    AXI_CLOCK_1_TO_0  = 8'd4,
    AXI_RESET_POSEDGE = 8'd5,
    AXI_RESET_NEGEDGE = 8'd6,
    AXI_RESET_ANYEDGE = 8'd7,
    AXI_RESET_0_TO_1  = 8'd8,
    AXI_RESET_1_TO_0  = 8'd9
} axi_wait_e;

`ifndef MAX_AXI_ADDRESS_WIDTH
  `define MAX_AXI_ADDRESS_WIDTH 64
`endif

`ifndef MAX_AXI_RDATA_WIDTH
  `define MAX_AXI_RDATA_WIDTH 1024
`endif

`ifndef MAX_AXI_WDATA_WIDTH
  `define MAX_AXI_WDATA_WIDTH 1024
`endif

`ifndef MAX_AXI_ID_WIDTH
  `define MAX_AXI_ID_WIDTH 18
`endif

// enum: axi_operation_mode_e
//
typedef enum int
{
    AXI_TRANSACTION_NON_BLOCKING = 32'd0,
    AXI_TRANSACTION_BLOCKING     = 32'd1
} axi_operation_mode_e;

// enum: axi_delay_mode_e
//
typedef enum int
{
    AXI_VALID2READY = 32'd0,
    AXI_TRANS2READY = 32'd1
} axi_delay_mode_e;

// enum: axi_write_data_mode_e
//
typedef enum int
{
    AXI_DATA_AFTER_ADDRESS = 32'd0,
    AXI_DATA_WITH_ADDRESS  = 32'd1
} axi_write_data_mode_e;

// Global Transaction Class
class axi_transaction;
    // Protocol 
    bit [((`MAX_AXI_ADDRESS_WIDTH) - 1):0]  addr;
    axi_size_e size;
    axi_burst_e burst;
    axi_lock_e lock;
    axi_cache_e cache;
    axi_prot_e prot;
    bit [((`MAX_AXI_ID_WIDTH) - 1):0]  id;
    bit [3:0] burst_length;
    bit [((((`MAX_AXI_RDATA_WIDTH > `MAX_AXI_WDATA_WIDTH) ? `MAX_AXI_RDATA_WIDTH : `MAX_AXI_WDATA_WIDTH)) - 1):0] data_words [];
    bit [(((`MAX_AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [];
    axi_response_e resp[];
    bit [7:0] addr_user;
    axi_rw_e read_or_write;
    int address_valid_delay;
    int data_valid_delay[];
    int write_response_valid_delay;
    int address_ready_delay;
    int data_ready_delay[];
    int write_response_ready_delay;

    // Housekeeping
    bit gen_write_strobes = 1'b1;
    axi_operation_mode_e  operation_mode  = AXI_TRANSACTION_BLOCKING;
    axi_delay_mode_e      delay_mode      = AXI_VALID2READY;
    axi_write_data_mode_e write_data_mode = AXI_DATA_WITH_ADDRESS;
    bit data_beat_done[];
    bit transaction_done;

    // This varaible is for printing component name and should not be visible/documented
    string driver_name;

    function void set_addr( input bit [((`MAX_AXI_ADDRESS_WIDTH) - 1):0]  laddr );
      addr = laddr;
    endfunction

    function bit [((`MAX_AXI_ADDRESS_WIDTH) - 1):0]   get_addr();
      return addr;
    endfunction

    function void set_size( input axi_size_e lsize );
      size = lsize;
    endfunction

    function axi_size_e get_size();
      return size;
    endfunction

    function void set_burst( input axi_burst_e lburst );
      burst = lburst;
    endfunction

    function axi_burst_e get_burst();
      return burst;
    endfunction

    function void set_lock( input axi_lock_e llock );
      lock = llock;
    endfunction

    function axi_lock_e get_lock();
      return lock;
    endfunction

    function void set_cache( input axi_cache_e lcache );
      cache = lcache;
    endfunction

    function axi_cache_e get_cache();
      return cache;
    endfunction

    function void set_prot( input axi_prot_e lprot );
      prot = lprot;
    endfunction

    function axi_prot_e get_prot();
      return prot;
    endfunction

    function void set_id( input bit [((`MAX_AXI_ID_WIDTH) - 1):0]  lid );
      id = lid;
    endfunction

    function bit [((`MAX_AXI_ID_WIDTH) - 1):0]   get_id();
      return id;
    endfunction

    function void set_burst_length( input bit [3:0] lburst_length );
      burst_length = lburst_length;
      data_words           = new[(lburst_length + 1)];
      write_strobes        = new[(lburst_length + 1)];
      resp                 = new[(lburst_length + 1)];
      data_valid_delay     = new[(lburst_length + 1)];
      data_ready_delay     = new[(lburst_length + 1)];
      data_beat_done       = new[(lburst_length + 1)];
    endfunction

    function bit [3:0]  get_burst_length();
      return burst_length;
    endfunction

    function void set_data_words( input bit [((((`MAX_AXI_RDATA_WIDTH > `MAX_AXI_WDATA_WIDTH) ? `MAX_AXI_RDATA_WIDTH : `MAX_AXI_WDATA_WIDTH)) - 1):0] ldata_words, input int index = 0 );
      data_words[index] = ldata_words;
    endfunction

    function bit [((((`MAX_AXI_RDATA_WIDTH > `MAX_AXI_WDATA_WIDTH) ? `MAX_AXI_RDATA_WIDTH : `MAX_AXI_WDATA_WIDTH)) - 1):0]  get_data_words( input int index = 0 );
      return data_words[index];
    endfunction

    function void set_write_strobes( input bit [(((`MAX_AXI_WDATA_WIDTH / 8)) - 1):0] lwrite_strobes, input int index = 0 );
      write_strobes[index] = lwrite_strobes;
    endfunction

    function bit [(((`MAX_AXI_WDATA_WIDTH / 8)) - 1):0]  get_write_strobes( input int index = 0 );
      return write_strobes[index];
    endfunction

    function void set_resp( input axi_response_e lresp, input int index = 0 );
      resp[index] = lresp;
    endfunction

    function axi_response_e get_resp( input int index = 0 );
      return resp[index];
    endfunction

    function void set_addr_user( input bit [7:0] laddr_user );
      addr_user = laddr_user;
    endfunction

    function bit [7:0]  get_addr_user();
      return addr_user;
    endfunction

    function void set_read_or_write( input axi_rw_e lread_or_write );
      read_or_write = lread_or_write;
    endfunction

    function axi_rw_e get_read_or_write();
      return read_or_write;
    endfunction

    function void set_address_valid_delay( input int laddress_valid_delay );
      address_valid_delay = laddress_valid_delay;
    endfunction

    function int get_address_valid_delay();
      return address_valid_delay;
    endfunction

    function void set_data_valid_delay( input int ldata_valid_delay, input int index = 0 );
      data_valid_delay[index] = ldata_valid_delay;
    endfunction

    function int get_data_valid_delay( input int index = 0 );
      return data_valid_delay[index];
    endfunction

    function void set_write_response_valid_delay( input int lwrite_response_valid_delay );
      write_response_valid_delay = lwrite_response_valid_delay;
    endfunction

    function int get_write_response_valid_delay();
      return write_response_valid_delay;
    endfunction

    function void set_address_ready_delay( input int laddress_ready_delay );
      address_ready_delay = laddress_ready_delay;
    endfunction

    function int get_address_ready_delay();
      return address_ready_delay;
    endfunction

    function void set_data_ready_delay( input int ldata_ready_delay, input int index = 0 );
      data_ready_delay[index] = ldata_ready_delay;
    endfunction

    function int get_data_ready_delay( input int index = 0 );
      return data_ready_delay[index];
    endfunction

    function void set_write_response_ready_delay( input int lwrite_response_ready_delay );
      write_response_ready_delay = lwrite_response_ready_delay;
    endfunction

    function int get_write_response_ready_delay();
      return write_response_ready_delay;
    endfunction

    function void set_gen_write_strobes( input bit lgen_write_strobes);
      gen_write_strobes = lgen_write_strobes;
    endfunction

    function bit get_gen_write_strobes();
      return gen_write_strobes;
    endfunction

    function void set_operation_mode( input axi_operation_mode_e loperation_mode );
      operation_mode = loperation_mode;
    endfunction

    function axi_operation_mode_e get_operation_mode();
      return operation_mode;
    endfunction

    function void set_delay_mode( input axi_delay_mode_e ldelay_mode );
      delay_mode = ldelay_mode;
    endfunction

    function axi_delay_mode_e get_delay_mode();
      return delay_mode;
    endfunction

    function void set_write_data_mode( input axi_write_data_mode_e lwrite_data_mode );
      write_data_mode = lwrite_data_mode;
    endfunction

    function axi_write_data_mode_e get_write_data_mode();
      return write_data_mode;
    endfunction

    function void set_data_beat_done( input int ldata_beat_done, input int index = 0 );
      data_beat_done[index] = ldata_beat_done;
    endfunction

    function int get_data_beat_done( input int index = 0 );
      return data_beat_done[index];
    endfunction

    function void set_transaction_done( input int ltransaction_done );
      transaction_done = ltransaction_done;
    endfunction

    function int get_transaction_done();
      return transaction_done;
    endfunction

    // Function: do_print
    //
    // Prints axi_transaction transaction attributes
    function void print (bit print_delays = 1'b0);
      $display("------------------------------------------------------------------------");
      $display("%0t: %s axi_transaction", $time, driver_name);
      $display("------------------------------------------------------------------------");
      $display("addr : 'h%h", addr);
      $display("size : %s", size.name());
      $display("burst : %s", burst.name());
      $display("lock : %s", lock.name());
      $display("cache : %s", cache.name());
      $display("prot : %s", prot.name());
      $display("id : 'h%h", id);
      $display("burst_length : 'h%h", burst_length);
      foreach( data_words[i0_1] )
        $display("data_words[%0d] : 'h%h", i0_1, data_words[i0_1]);
      foreach( write_strobes[i0_1] )
        $display("write_strobes[%0d] : 'h%h", i0_1, write_strobes[i0_1]);
      foreach( resp[i0_1] )
        $display("resp[%0d] : %s", i0_1, resp[i0_1].name());
      $display("addr_user : 'h%h", addr_user);
      $display("read_or_write : %s", read_or_write.name());
      $display("gen_write_strobes : 'b%b", gen_write_strobes );
      $display("operation_mode   : %s", operation_mode.name() );
      $display("delay_mode       : %s", delay_mode.name() );
      $display("write_data_mode  : %s", write_data_mode.name() );
      foreach( data_beat_done[i0_1] )
        $display("data_beat_done[%0d] : 'b%b", i0_1, data_beat_done[i0_1] );
      $display("transaction_done : 'b%b", transaction_done );
      if ( print_delays == 1'b1 )
      begin
        $display("address_valid_delay : %0d", address_valid_delay);
        foreach( data_valid_delay[i0_1] )
          $display("data_valid_delay[%0d] : %0d", i0_1, data_valid_delay[i0_1]);
        $display("write_response_valid_delay : %0d", write_response_valid_delay);
        $display("address_ready_delay : %0d", address_ready_delay);
        foreach( data_ready_delay[i0_1] )
          $display("data_ready_delay[%0d] : %0d", i0_1, data_ready_delay[i0_1]);
        $display("write_response_ready_delay : %0d", write_response_ready_delay);
      end
    endfunction
endclass

`else
// *****************************************************************************
//
// Copyright 2007-2016 Mentor Graphics Corporation
// All Rights Reserved.
//
// THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE PROPERTY OF
// MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS.
//
// *****************************************************************************
// SystemVerilog           Version: 20160107
// *****************************************************************************

// Title: AXI Enumeration Types
//

//------------------------------------------------------------------------------
//
// Enum: axi_size_e
//
//------------------------------------------------------------------------------
//  Word size encoding 
typedef enum bit [2:0]
{
    AXI_BYTES_1   = 3'h0,
    AXI_BYTES_2   = 3'h1,
    AXI_BYTES_4   = 3'h2,
    AXI_BYTES_8   = 3'h3,
    AXI_BYTES_16  = 3'h4,
    AXI_BYTES_32  = 3'h5,
    AXI_BYTES_64  = 3'h6,
    AXI_BYTES_128 = 3'h7
} axi_size_e;



//------------------------------------------------------------------------------
//
// Enum: axi_prot_e
//
//------------------------------------------------------------------------------
//  Protection type 
typedef enum bit [2:0]
{
    AXI_NORM_SEC_DATA    = 3'h0,
    AXI_PRIV_SEC_DATA    = 3'h1,
    AXI_NORM_NONSEC_DATA = 3'h2,
    AXI_PRIV_NONSEC_DATA = 3'h3,
    AXI_NORM_SEC_INST    = 3'h4,
    AXI_PRIV_SEC_INST    = 3'h5,
    AXI_NORM_NONSEC_INST = 3'h6,
    AXI_PRIV_NONSEC_INST = 3'h7
} axi_prot_e;



//------------------------------------------------------------------------------
//
// Enum: axi_cache_e
//
//------------------------------------------------------------------------------
//  Cache type
typedef enum bit [3:0]
{
    AXI_NONCACHE_NONBUF             = 4'h0,
    AXI_BUF_ONLY                    = 4'h1,
    AXI_CACHE_NOALLOC               = 4'h2,
    AXI_CACHE_BUF_NOALLOC           = 4'h3,
    AXI_CACHE_RSVD0                 = 4'h4,
    AXI_CACHE_RSVD1                 = 4'h5,
    AXI_CACHE_WTHROUGH_ALLOC_R_ONLY = 4'h6,
    AXI_CACHE_WBACK_ALLOC_R_ONLY    = 4'h7,
    AXI_CACHE_RSVD2                 = 4'h8,
    AXI_CACHE_RSVD3                 = 4'h9,
    AXI_CACHE_WTHROUGH_ALLOC_W_ONLY = 4'ha,
    AXI_CACHE_WBACK_ALLOC_W_ONLY    = 4'hb,
    AXI_CACHE_RSVD4                 = 4'hc,
    AXI_CACHE_RSVD5                 = 4'hd,
    AXI_CACHE_WTHROUGH_ALLOC_RW     = 4'he,
    AXI_CACHE_WBACK_ALLOC_RW        = 4'hf
} axi_cache_e;



//------------------------------------------------------------------------------
//
// Enum: axi_burst_e
//
//------------------------------------------------------------------------------
//  This specifies Burst type which determines address calculation
typedef enum bit [1:0]
{
    AXI_FIXED      = 2'h0,
    AXI_INCR       = 2'h1,
    AXI_WRAP       = 2'h2,
    AXI_BURST_RSVD = 2'h3
} axi_burst_e;



//------------------------------------------------------------------------------
//
// Enum: axi_response_e
//
//------------------------------------------------------------------------------
//  Response type 
typedef enum bit [1:0]
{
    AXI_OKAY   = 2'h0,
    AXI_EXOKAY = 2'h1,
    AXI_SLVERR = 2'h2,
    AXI_DECERR = 2'h3
} axi_response_e;



//------------------------------------------------------------------------------
//
// Enum: axi_lock_e
//
//------------------------------------------------------------------------------
//  Lock type for atomic accesses
typedef enum bit [1:0]
{
    AXI_NORMAL    = 2'h0,
    AXI_EXCLUSIVE = 2'h1,
    AXI_LOCKED    = 2'h2,
    AXI_LOCK_RSVD = 2'h3
} axi_lock_e;



//------------------------------------------------------------------------------
//
// Enum: axi_rw_e
//
//------------------------------------------------------------------------------
//  Specifies transaction type read or write 
typedef enum bit [0:0]
{
    AXI_TRANS_READ  = 1'h0,
    AXI_TRANS_WRITE = 1'h1
} axi_rw_e;



//------------------------------------------------------------------------------
//
// Enum: axi_len_e
//
//------------------------------------------------------------------------------
//  Specifies length of the transaction 
typedef enum bit [3:0]
{
    AXI_LENGTH_1  = 4'h0,
    AXI_LENGTH_2  = 4'h1,
    AXI_LENGTH_3  = 4'h2,
    AXI_LENGTH_4  = 4'h3,
    AXI_LENGTH_5  = 4'h4,
    AXI_LENGTH_6  = 4'h5,
    AXI_LENGTH_7  = 4'h6,
    AXI_LENGTH_8  = 4'h7,
    AXI_LENGTH_9  = 4'h8,
    AXI_LENGTH_10 = 4'h9,
    AXI_LENGTH_11 = 4'ha,
    AXI_LENGTH_12 = 4'hb,
    AXI_LENGTH_13 = 4'hc,
    AXI_LENGTH_14 = 4'hd,
    AXI_LENGTH_15 = 4'he,
    AXI_LENGTH_16 = 4'hf
} axi_len_e;



//------------------------------------------------------------------------------
//
// Enum: axi_error_e
//
//------------------------------------------------------------------------------
//  Specifies error type 
typedef enum bit [3:0]
{
    AXI_AWBURST_RSVD        = 4'h0,
    AXI_ARBURST_RSVD        = 4'h1,
    AXI_AWSIZE_GT_BUS_WIDTH = 4'h2,
    AXI_ARSIZE_GT_BUS_WIDTH = 4'h3,
    AXI_AWLOCK_RSVD         = 4'h4,
    AXI_ARLOCK_RSVD         = 4'h5,
    AXI_AWLEN_LAST_MISMATCH = 4'h6,
    AXI_AWID_WID_MISMATCH   = 4'h7,
    AXI_WSTRB_ILLEGAL       = 4'h8,
    AXI_AWCACHE_RSVD        = 4'h9,
    AXI_ARCACHE_RSVD        = 4'ha
} axi_error_e;



//------------------------------------------------------------------------------
//
// Enum: axi_assertion_e
//
//------------------------------------------------------------------------------
//  Type defining the assertion messages which can be produced by the <mgc_axi> QVIP.
// 
// Individual assertion messages can be disabled using the <config_enable_assertion> array of configuration bits.
// 
// AXI_ARESETn_SIGNAL_Z                                                        -  60000 -  AXI reset signal (ARESETn) has a value Z
// AXI_ARESETn_SIGNAL_X                                                        -  60001 -  AXI reset signal (ARESETn) has a value X
// AXI_ACLK_SIGNAL_Z                                                           -  60002 -  
// AXI_ADDR_FOR_READ_BURST_ACROSS_4K_BOUNDARY                                  -  60004 -  This read transaction has crossed a 4KB boundary (SPEC3(A3.4.1))
// AXI_ADDR_FOR_WRITE_BURST_ACROSS_4K_BOUNDARY                                 -  60005 -  This write transaction has crossed a 4KB boundary (SPEC3(A3.4.1))
// AXI_ARADDR_CHANGED_BEFORE_ARREADY                                           -  60006 -  The value of <ARADDR> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARADDR_UNKN                                                             -  60007 -  <ARADDR> has an X value/<ARADDR> has an Z value (SPEC3(A2.5))
// AXI_ARBURST_CHANGED_BEFORE_ARREADY                                          -  60008 -  The value of <ARBURST> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARBURST_UNKN                                                            -  60009 -  <ARBURST> has an X value/<ARBURST> has an Z value (SPEC3(A2.5))
// AXI_ARCACHE_CHANGED_BEFORE_ARREADY                                          -  60010 -  The value of <ARCACHE> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARCACHE_UNKN                                                            -  60011 -  <ARCACHE> has an X value/<ARCACHE> has an Z value (SPEC3(A2.5))
// AXI_ARID_CHANGED_BEFORE_ARREADY                                             -  60012 -  The value of <ARID> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARID_UNKN                                                               -  60013 -  <ARID> has an X value/<ARID> has an Z value (SPEC3(A2.5))
// AXI_ARLEN_CHANGED_BEFORE_ARREADY                                            -  60014 -  The value of <ARLEN> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARLEN_UNKN                                                              -  60015 -  <ARLEN> has an X value/<ARLEN> has an Z value (SPEC3(A2.5))
// AXI_ARLOCK_CHANGED_BEFORE_ARREADY                                           -  60016 -  The value of <ARLOCK> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARLOCK_UNKN                                                             -  60017 -  <ARLOCK> has an X value/<ARLOCK> has an Z value (SPEC3(A2.5))
// AXI_ARPROT_CHANGED_BEFORE_ARREADY                                           -  60018 -  The value of <ARPROT> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARPROT_UNKN                                                             -  60019 -  <ARPROT> has an X value/<ARPROT> has an Z value (SPEC3(A2.5))
// AXI_ARREADY_UNKN                                                            -  60020 -  <ARREADY> has an X value/<ARREADY> has a Z value (SPEC3(A2.5))
// AXI_ARSIZE_CHANGED_BEFORE_ARREADY                                           -  60021 -  The value of <ARSIZE> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARSIZE_UNKN                                                             -  60022 -  <ARSIZE> has an X value/<ARSIZE> has an Z value (SPEC3(A2.5))
// AXI_ARUSER_CHANGED_BEFORE_ARREADY                                           -  60023 -  The value of <ARUSER> has changed from its initial value between the time <ARVALID> was asserted, and before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARUSER_UNKN                                                             -  60024 -  <ARUSER> has an X value/<ARUSER> has an Z value (SPEC3(A2.5))
// AXI_ARVALID_DEASSERTED_BEFORE_ARREADY                                       -  60025 -  <ARVALID> has been de-asserted before <ARREADY> was asserted (SPEC3(A3.2.1))
// AXI_ARVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                 -  60026 -  A master interface must begin driving <ARVALID> high only at a rising clock edge after <ARESETn> is HIGH (SPEC3(A3.1.2))
// AXI_ARVALID_UNKN                                                            -  60027 -  <ARVALID> has an X value/<ARVALID> has an Z value (SPEC3(A2.5))
// AXI_AWADDR_CHANGED_BEFORE_AWREADY                                           -  60028 -  The value of <AWADDR> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))
// AXI_AWADDR_UNKN                                                             -  60029 -  <AWADDR> has an X value/<AWADDR> has an Z value (SPEC3(A2.2))
// AXI_AWBURST_CHANGED_BEFORE_AWREADY                                          -  60030 -  The value of <AWBURST> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))
// AXI_AWBURST_UNKN                                                            -  60031 -  <AWBURST> has an X value/<AWBURST> has an Z value (SPEC3(A2.2))
// AXI_AWCACHE_CHANGED_BEFORE_AWREADY                                          -  60032 -  The value of <AWCACHE> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                       
// AXI_AWCACHE_UNKN                                                            -  60033 -  <AWCACHE> has an X value/AWCACHE has an Z value (SPEC3(A2.2))
// AXI_AWID_CHANGED_BEFORE_AWREADY                                             -  60034 -  The value of <AWID> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))
// AXI_AWID_UNKN                                                               -  60035 -  <AWID> has an X value/<AWID> has an Z value (SPEC3(A2.2))
// AXI_AWLEN_CHANGED_BEFORE_AWREADY                                            -  60036 -  The value of <AWLEN> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))
// AXI_AWLEN_UNKN                                                              -  60037 -  <AWLEN> has an X value/<AWLEN> has an Z value (SPEC3(A2.2))                                                                                                                                        
// AXI_AWLOCK_CHANGED_BEFORE_AWREADY                                           -  60038 -  The value of <AWLOCK> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                            
// AXI_AWLOCK_UNKN                                                             -  60039 -  <AWLOCK> has an X value/<AWLOCK> has an Z value (SPEC3(A2.2))
// AXI_AWPROT_CHANGED_BEFORE_AWREADY                                           -  60040 -  The value of <AWPROT> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                          
// AXI_AWPROT_UNKN                                                             -  60041 -  <AWPROT> has an X value/<AWPROT> has an Z value (SPEC3(A2.2))                                                                                                                                        
// AXI_AWREADY_UNKN                                                            -  60042 -  <AWREADY> has an X value/<AWREADY> has an Z value (SPEC3(A2.2))                                                                                                                                        
// AXI_AWSIZE_CHANGED_BEFORE_AWREADY                                           -  60043 -  The value of <AWSIZE> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                                       
// AXI_AWSIZE_UNKN                                                             -  60044 -  <AWSIZE> has an X value/<AWSIZE> has an Z value (SPEC3(A2.2))                                                                                                                                                 
// AXI_AWUSER_CHANGED_BEFORE_AWREADY                                           -  60045 -  The value of <AWUSER> has changed from its initial value between the time <AWVALID> was asserted, and before <AWREADY> was asserted (SPEC3(A3.2.1))                                           
// AXI_AWUSER_UNKN                                                             -  60046 -  <AWUSER> has an X value/<AWUSER> has an Z value (SPEC3(A3.1))                                                                                                                                                    
// AXI_AWVALID_DEASSERTED_BEFORE_AWREADY                                       -  60047 -  <AWVALID> has been de-asserted before <AWREADY> was asserted (SPEC3(A3.2.2))                                                                                                                  
// AXI_AWVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                 -  60048 -  A master interface must begin driving <AWVALID> high only at a rising clock edge after <ARESETn> is HIGH (SPEC3(A3.1.2))                                                               
// AXI_AWVALID_UNKN                                                            -  60049 -  <AWVALID> has an X value/<AWVALID> has an Z value (SPEC3(A2.2))                                                                                                                                                 
// AXI_BID_CHANGED_BEFORE_BREADY                                               -  60050 -  The value of <BID> has changed from its initial value between the time <BVALID> was asserted, and before <BREADY> was asserted (SPEC3(A3.2.1))                                                 
// AXI_BID_UNKN                                                                -  60051 -  <BID> has an X value/<BID> has a Z value (SPEC3(A2.4))                                                                                                                                                       
// AXI_BREADY_UNKN                                                             -  60052 -  <BREADY> has an X value/<BREADY> has an Z value (SPEC3(A2.4))                                                                                                                                                 
// AXI_BRESP_CHANGED_BEFORE_BREADY                                             -  60053 -  The value of <BRESP> has changed from its initial value between the time <BVALID> was asserted, and before <BREADY> was asserted (SPEC3(A3.2.1))                                            
// AXI_BRESP_UNKN                                                              -  60054 -  <BRESP> has an X value/<BRESP> has a Z value (SPEC3(A2.4))                                                                                                                                                   
// AXI_BUSER_CHANGED_BEFORE_BREADY                                             -  60055 -  The value of <BUSER> has changed from its initial value between the time <BVALID> was asserted, and before <BREADY> was asserted (SPEC3(A3.2.1))                                       
// AXI_BUSER_UNKN                                                              -  60056 -  <BUSER> has an X value/<BUSER> has a Z value (SPEC3(A2.4))                                                                                                                                                       
// AXI_BVALID_DEASSERTED_BEFORE_BREADY                                         -  60057 -  <BVALID> has been de-asserted before <BREADY> was asserted (SPEC3(A3.2.1))                                                                                                                       
// AXI_BVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  -  60058 -  A slave interface must begin driving  <BVALID> high only at a rising clock edge after ARESETn is HIGH (SPEC3(A3.1.2))                                                                        
// AXI_BVALID_UNKN                                                             -  60059 -  <BVALID> has an X value/<BVALID> has a Z value (SPEC3(A2.4))                                                                                                                                                   
// AXI_EXCLUSIVE_READ_ACCESS_MODIFIABLE                                        -  60060 -  The modifiable bit (bit 1 of the cache parameter) should not be set for an exclusive read access (SPEC3(A7.2.4))                                                                                 
// AXI_EXCLUSIVE_READ_BYTES_TRANSFER_EXCEEDS_128                               -  60061 -  Number of bytes in an exclusive read transaction must be less than or equal to 128 (SPEC3(A7.2.4))                                                                                         
// AXI_EXCLUSIVE_WRITE_BYTES_TRANSFER_EXCEEDS_128                              -  60062 -  Number of bytes in an exclusive write transaction must be less than or equal to 128 (SPEC3(A7.2.4))                                                                                
// AXI_EXCLUSIVE_READ_BYTES_TRANSFER_NOT_POWER_OF_2                            -  60063 -  Number of bytes of an exclusive read transaction is not a power of 2 (SPEC3(A7.2.4))                                                                                           
// AXI_EXCLUSIVE_WRITE_BYTES_TRANSFER_NOT_POWER_OF_2                           -  60064 -  Number of bytes of an exclusive write transaction is not a power of 2 (SPEC3(A7.2.4))                                                                                               
// AXI_EXCLUSIVE_WR_ADDRESS_NOT_SAME_AS_RD                                     -  60065 -  Exclusive write does not match the address of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                                        
// AXI_EXCLUSIVE_WR_BURST_NOT_SAME_AS_RD                                       -  60066 -  Exclusive write does not match the burst setting of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                                      
// AXI_EXCLUSIVE_WR_CACHE_NOT_SAME_AS_RD                                       -  60067 -  Exclusive write does not match the cache setting of the previous exclusive read to this id (see the ARM AXI compliance-checker AXI_RECM_EXCL_MATCH assertion code) (SPEC3(A7.2.4))            
// AXI_EXCLUSIVE_WRITE_ACCESS_MODIFIABLE                                       -  60068 -  The modifiable bit (bit 1 of the cache parameter) should not be set for an exclusive write access (SPEC3(A7.2.4))                                                               
// AXI_EXCLUSIVE_WR_LENGTH_NOT_SAME_AS_RD                                      -  60069 -  Exclusive write does not match the length of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                           
// AXI_EXCLUSIVE_WR_PROT_NOT_SAME_AS_RD                                        -  60070 -  Exclusive write does not match the prot setting of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                       
// AXI_EXCLUSIVE_WR_SIZE_NOT_SAME_AS_RD                                        -  60071 -  Exclusive write does not match the size of the previous exclusive read to this id (SPEC3(A7.2.4))                                                                               
// AXI_EXOKAY_RESPONSE_NORMAL_READ                                             -  60072 -  Slave has responded ~AXI_EXOKAY~ to a non exclusive read transfer                                                                                                                
// AXI_EXOKAY_RESPONSE_NORMAL_WRITE                                            -  60073 -  Slave has responded ~AXI_EXOKAY~ to a non exclusive write transfer                                                                                                               
// AXI_EX_RD_RESP_MISMATCHED_WITH_EXPECTED_RESP                                -  60074 -  Expected response to this exclusive read did not matched with the actual response (SPEC3(A7.2.3))                                                                            
// AXI_EX_WR_RESP_MISMATCHED_WITH_EXPECTED_RESP                                -  60075 -  Expected response to this exclusive write did not matched with the actual response (SPEC3(A7.2.3))                                                                           
// AXI_EX_RD_EXOKAY_RESP_SLAVE_WITHOUT_EXCLUSIVE_ACCESS                        -  60076 -  Response for an exclusive read to a slave which does not support exclusive access should be ~AXI_OKAY~, but it returned ~AXI_EXOKAY~ (SPEC3(A7.2.3))
// AXI_EX_WRITE_BEFORE_EX_READ_RESPONSE                                        -  60077 -  Exclusive write has occurred, with no previous exclusive read (SPEC3(A7.2.2))                                                                                                        
// AXI_EX_WRITE_EXOKAY_RESP_SLAVE_WITHOUT_EXCLUSIVE_ACCESS                     -  60078 -  Response for an exclusive write to a slave which does not support exclusive access should be ~AXI_OKAY~, but it returned ~AXI_EXOKAY~ (SPEC3(A7.2.3))              
// AXI_ILLEGAL_LENGTH_WRAPPING_READ_BURST                                      -  60079 -  In the last read address phase burst_length has an illegal value for a burst of type AXI_WRAP (SPEC3(A3.4.1))                                                         
// AXI_ILLEGAL_LENGTH_WRAPPING_WRITE_BURST                                     -  60080 -  In the last write address phase burst_length has an illegal value for a burst of type AXI_WRAP (SPEC3(A3.4.1))                                                        
// AXI_ILLEGAL_RESPONSE_EXCLUSIVE_READ                                         -  60081 -  Response for an exclusive read should be either ~AXI_OKAY~ or ~AXI_EXOKAY~ (SPEC3(A7.2.3))                                                                                    
// AXI_ILLEGAL_RESPONSE_EXCLUSIVE_WRITE                                        -  60082 -  Response for an exclusive write should be either ~AXI_OKAY~ or ~AXI_EXOKAY~ (SPEC3(A7.2.3))                                                                                   
// AXI_PARAM_READ_DATA_BUS_WIDTH                                               -  60083 -  The value of <AXI_RDATA_WIDTH> must be one of 8,16,32,64,128,256,512,1024 (SPEC3(A1.3.1))                                                                                            
// AXI_PARAM_WRITE_DATA_BUS_WIDTH                                              -  60084 -  The value of <AXI_WDATA_WIDTH> must be one of 8,16,32,64,128,256,512,1024 (SPEC3(A1.3.1))                                                                                        
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_12                                    -  60085 -  The RA bit of the cache parameter should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                              
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_13                                    -  60086 -  The RA bit of the cache parameter should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                             
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_4                                     -  60087 -  The RA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                                
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_5                                     -  60088 -  The RA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                                  
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_8                                     -  60089 -  The RA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                                     
// AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_9                                     -  60090 -  The RA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                                                                     
// AXI_READ_BURST_LENGTH_VIOLATION                                             -  60091 -  The burst_length implied by the number of beats actually read does not match the burst_length defined by the <axi_master_read_addr_channel_phase> (SPEC3(A3.4.1))                             
// AXI_READ_BURST_SIZE_VIOLATION                                               -  60092 -  In this read transaction, size has been set greater than the defined data bus width (SPEC3(A3.4.1))                                                                                                   
// AXI_READ_DATA_BEFORE_ADDRESS                                                -  60093 -  An unexpected read response has occurred (there are no outstanding read transactions with this id) (SPEC3(A3.3.1))                                                                           
// AXI_READ_DATA_CHANGED_BEFORE_RREADY                                         -  60094 -  The value of <RDATA> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                              
// AXI_READ_DATA_UNKN                                                          -  60095 -  <RDATA> has an X value/<RDATA> has a Z value (SPEC3(A2.6))                                                                                                                                     
// AXI_RESERVED_ARLOCK_ENCODING                                                -  60096 -  The reserved encoding of 2'b11 should not be used for ARLOCK (SPEC3(A7.4))                                                                                                                   
// AXI_READ_RESP_CHANGED_BEFORE_RREADY                                         -  60097 -  The value of <RRESP> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                        
// AXI_RESERVED_ARBURST_ENCODING                                               -  60098 -  The reserved encoding of 2'b11 should not be used for <ARBURST> (SPEC3(A3.4.1))                                                                                              
// AXI_RESERVED_AWBURST_ENCODING                                               -  60099 -  The reserved encoding of 2'b11 should not be used for <AWBURST> (SPEC3(A3.4.1))                                                                                                  
// AXI_RID_CHANGED_BEFORE_RREADY                                               -  60100 -  The value of <RID> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                              
// AXI_RID_UNKN                                                                -  60101 -  <RID> has an X value/<RID> has a Z value (SPEC3(A2.6))                                                                                                                                    
// AXI_RLAST_CHANGED_BEFORE_RREADY                                             -  60102 -  The value of <RLAST> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                     
// AXI_RLAST_UNKN                                                              -  60103 -  <RLAST> has an X value/<RLAST> has a Z value (SPEC3(A2.6))                                                                                                                                 
// AXI_RREADY_UNKN                                                             -  60104 -  <RREADY> has an X value/<RREADY> has a Z value (SPEC3(A2.6))                                                                                                                                   
// AXI_RRESP_UNKN                                                              -  60105 -  <RRESP> has an X value/<RRESP> has a Z value (SPEC3(A2.6))                                                                                                                                  
// AXI_RUSER_CHANGED_BEFORE_RREADY                                             -  60106 -  The value of <RUSER> has changed from its initial value between the time <RVALID> was asserted, and before <RREADY> was asserted (SPEC3(A3.2.1))                          
// AXI_RUSER_UNKN                                                              -  60107 -  <RUSER> has an X value/<RUSER> has a Z value (SPEC3(A2.6))                                                                                                              
// AXI_RVALID_DEASSERTED_BEFORE_RREADY                                         -  60108 -  <RVALID> has been de-asserted before <RREADY> was asserted (SPEC3(A3.2.1))                                                                         
// AXI_RVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  -  60109 -  A slave interface must begin driving  <RVALID> high only at a rising clock edge after ARESETn is HIGH (SPEC3(A3.1.2))                                  
// AXI_RVALID_UNKN                                                             -  60110 -  <RVALID> has an X value/<RVALID> has a Z value (SPEC3(A2.6))                                                                                                        
// AXI_UNALIGNED_ADDRESS_FOR_EXCLUSIVE_READ                                    -  60111 -  Exclusive read accesses must have address aligned to the total number of bytes in the transaction (SPEC3(A7.2.4))                                     
// AXI_UNALIGNED_ADDRESS_FOR_EXCLUSIVE_WRITE                                   -  60112 -  Exclusive write accesses must have address aligned to the total number of bytes in the transaction (SPEC3(A7.2.4))                                     
// AXI_UNALIGNED_ADDR_FOR_WRAPPING_READ_BURST                                  -  60113 -  Wrapping bursts must have address aligned to the start of the read transfer (SPEC3(A3.4.1))                                                                                                                                    
// AXI_UNALIGNED_ADDR_FOR_WRAPPING_WRITE_BURST                                 -  60114 -  Wrapping bursts must have address aligned to the start of the write transfet (SPEC3(A3.4.1))                                                                                                                                    
// AXI_WDATA_CHANGED_BEFORE_WREADY_ON_INVALID_LANE                             -  60115 -  On a lane whose strobe is 0, the value of <WDATA> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                               
// AXI_WDATA_CHANGED_BEFORE_WREADY_ON_VALID_LANE                               -  60116 -  On a lane whose strobe is 1, the value of <WDATA> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                   
// AXI_WLAST_CHANGED_BEFORE_WREADY                                             -  60117 -  The value of <WLAST> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                
// AXI_WID_CHANGED_BEFORE_WREADY                                               -  60118 -  The value of <WID> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                
// AXI_WLAST_UNKN                                                              -  60119 -  <WLAST> has an X value/<WLAST> has an Z value (SPEC3(A2.3))                                                                                        
// AXI_WID_UNKN                                                                -  60120 -  <WID> has an X value/<WID> has an Z value (SPEC3(A2.3))                                                                                                     
// AXI_WREADY_UNKN                                                             -  60121 -  <WREADY> has an X value/<WREADY> has a Z value (SPEC3(A2.3))                                                                                       
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_12                                   -  60122 -  The WA bit of the cache parameter should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                     
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_13                                   -  60123 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                   
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_4                                    -  60124 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                              
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_5                                    -  60125 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                         
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_8                                    -  60126 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                           
// AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_9                                    -  60127 -  The WA of the cache parameter bit should not be HIGH when the Modifiable bit is LOW (SPEC3(A4.4))                                            
// AXI_WRITE_BURST_SIZE_VIOLATION                                              -  60128 -  In this write transaction, size has been set greater than the defined data buswidth (SPEC3(A3.4.1))                                         
// AXI_WRITE_DATA_BEFORE_ADDRESS                                               -  60129 -  A write data beat has occurred before the corresponding address phase                                                                      
// AXI_WRITE_DATA_UNKN_ON_INVALID_LANE                                         -  60130 -  DEPRECATED - This assertion is now DEPRECATED and by default DISABLED, as per protocol Byte lanes for which strobe is 0 could take unknown value..
// AXI_WRITE_DATA_UNKN_ON_VALID_LANE                                           -  60131 -  On a lane whose strobe is 1, <WDATA> has an X value/<WDATA> has a Z value (SPEC3(A2.3))                                          
// AXI_RESERVED_AWLOCK_ENCODING                                                -  60132 -  The reserved encoding of 2'b11 should not be used for AWLOCK (SPEC3(A7.4))                                                                                                                                
// AXI_WRITE_STROBE_ON_INVALID_BYTE_LANES                                      -  60133 -  Write strobe(s) incorrect for the address/size of a fixed transfer (SPEC3(A2.3))                                                                                                                  
// AXI_WSTRB_CHANGED_BEFORE_WREADY                                             -  60134 -  The value of <WSTRB> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                         
// AXI_WSTRB_UNKN                                                              -  60135 -  <WSTRB> has an X value/<WSTRB> has an Z value (SPEC3(A2.3))                                                                                                                                                      
// AXI_WUSER_CHANGED_BEFORE_WREADY                                             -  60136 -  The value of <WUSER> has changed from its initial value between the time <WVALID> was asserted, and before <WREADY> was asserted (SPEC3(A3.2.1))                                        
// AXI_WUSER_UNKN                                                              -  60137 -  <WUSER> has an X value/<WUSER> has an Z value (SPEC3(A2.3))                                                                                                                              
// AXI_WVALID_DEASSERTED_BEFORE_WREADY                                         -  60138 -  <WVALID> has been de-asserted before <WREADY> was asserted (SPEC3(A3.2.1))                                                                                               
// AXI_WVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  -  60139 -  A master interface must begin driving <WVALID> high only at a rising clock edge after <ARESETn> is HIGH (SPEC3(A3.1.2))                                             
// AXI_WVALID_UNKN                                                             -  60140 -  <WVALID> has an X value/<WVALID> has an Z value (SPEC3(A2.3))                                                                                                             
// AXI_ADDR_ACROSS_4K_WITHIN_LOCKED_WRITE_TRANSACTION                          -  60141 -  Transactions within a locked write sequence should be within the same 4K address boundary (SPEC3(A7.3))                                           
// AXI_ADDR_ACROSS_4K_WITHIN_LOCKED_READ_TRANSACTION                           -  60142 -  Transactions within a locked read sequence should be within the same 4K address boundary (SPEC3(A7.3))                                            
// AXI_AWID_CHANGED_WITHIN_LOCKED_TRANSACTION                                  -  60143 -  Master should not change the awid within the locked transaction (SPEC3(A7.3))                                               
// AXI_ARID_CHANGED_WITHIN_LOCKED_TRANSACTION                                  -  60144 -  Master should not change the arid within the locked transaction (SPEC3(A7.3))                                              
// AXI_AWPROT_CHANGED_WITHIN_LOCKED_TRANSACTION                                -  60145 -  Master should not change the awprot within the locked transaction (SPEC3(A7.3))                                                   
// AXI_ARPROT_CHANGED_WITHIN_LOCKED_TRANSACTION                                -  60146 -  Master should not change the arprot within the locked transaction (SPEC3(A7.3))                                                 
// AXI_AWCACHE_CHANGED_WITHIN_LOCKED_TRANSACTION                               -  60147 -  Master should not change the awcache within the locked transaction (SPEC3(A7.3))                                                    
// AXI_ARCACHE_CHANGED_WITHIN_LOCKED_TRANSACTION                               -  60148 -  Master should not change the arcache within the locked transaction (SPEC3(A7.3))                                                      
// AXI_NUMBER_OF_LOCKED_SEQUENCES_EXCEEDS_2                                    -  60149 -  Number of accesses within a locked sequence should not be more than 2 (SPEC3(A7.3))                                                                                                     
// AXI_LOCKED_WRITE_BEFORE_COMPLETION_OF_PREVIOUS_WRITE_TRANSACTIONS           -  60150 -  A locked write sequence should not commence before completion of all previously issued write addresses (SPEC3(A7.3))                                                 
// AXI_LOCKED_WRITE_BEFORE_COMPLETION_OF_PREVIOUS_READ_TRANSACTIONS            -  60151 -  A locked write sequence should not commence before completion of all previously issued read addresses (SPEC3(A7.3))                                              
// AXI_LOCKED_READ_BEFORE_COMPLETION_OF_PREVIOUS_WRITE_TRANSACTIONS            -  60152 -  A locked read sequence should not commence before completion of all previously issued write addresses (SPEC3(A7.3))                                                    
// AXI_LOCKED_READ_BEFORE_COMPLETION_OF_PREVIOUS_READ_TRANSACTIONS             -  60153 -  A locked read sequence should not commence before completion of all previously issued read addresses (SPEC3(A7.3))                                                        
// AXI_NEW_BURST_BEFORE_COMPLETION_OF_UNLOCK_TRANSACTION                       -  60154 -  The unlocking transaction should be completed before further any transactions are initiated (SPEC3(A7.3))                                                           
// AXI_UNLOCKED_WRITE_WHILE_OUTSTANDING_LOCKED_WRITES                          -  60155 -  Unlocking write transaction started while outstanding locked write transaction has not completed (SPEC3(A7.3))                                                  
// AXI_UNLOCKED_WRITE_WHILE_OUTSTANDING_LOCKED_READS                           -  60156 -  Unlocking write transaction started while outstanding locked read transaction has not completed (SPEC3(A7.3))                                                 
// AXI_UNLOCKED_READ_WHILE_OUTSTANDING_LOCKED_WRITES                           -  60157 -  Unlocking read transaction started while outstanding locked write transaction has not completed (SPEC3(A7.3))                                                             
// AXI_UNLOCKED_READ_WHILE_OUTSTANDING_LOCKED_READS                            -  60158 -  Unlocking read transaction started while outstanding locked read transaction has not completed (SPEC3(A7.3))                                                     
// AXI_UNLOCKING_TRANSACTION_WITH_AN_EXCLUSIVE_ACCESS                          -  60159 -  Unlocking transaction can not be an exclusive access transaction (SPEC3(A7.3))                                                                                                                                                            
// AXI_FIRST_DATA_ITEM_OF_TRANSACTION_WRITE_ORDER_VIOLATION                    -  60160 -  The order in which a slave receives the first data item of each transaction must be the same as the order in which it receives the addresses for the transaction (SPEC3(A5.3.3))                                                      
// AXI_AWLEN_MISMATCHED_WITH_COMPLETED_WRITE_DATA_BURST                        -  60161 -  AWLEN value of write address control does not match with corresponding outstanding write data burts length (SPEC3(A3.4.1))                                                       
// AXI_WRITE_LENGTH_MISMATCHED_ACTUAL_LENGTH_OF_WRITE_DATA_BURST_EXCEEDS_AWLEN -  60162 -  The actual length of write data burst exceeds with the length specified by AWLEN (SPEC3(A3.4.1))                                              
// AXI_AWLEN_MISMATCHED_ACTUAL_LENGTH_OF_WRITE_DATA_BURST_EXCEEDS_AWLEN        -  60163 -  Actual length of data burst has exceeded the burst length specified by AWLEN (SPEC3(A3.4.1))                                                               
// AXI_WLAST_ASSERTED_DURING_DATA_PHASE_OTHER_THAN_LAST                        -  60164 -  AWLEN value of write address control does not match with corresponding outstanding write data burts length (SPEC3(A3.4.1))                                                 
// AXI_WRITE_INTERLEAVE_DEPTH_VIOLATION                                        -  60165 -  Write data bursts should not be interleaved beyond the write interleaving depth (SPEC3(A5.3.3))                                   
// AXI_WRITE_RESPONSE_WITHOUT_ADDR                                             -  60166 -  Write response should not be sent before the corresponding address has completed (SPEC3(A3.3.1))                                 
// AXI_WRITE_RESPONSE_WITHOUT_DATA                                             -  60167 -  Write response should not be sent before the corresponding write data burst completed (SPEC3(A3.3.1))                           
// AXI_AWVALID_HIGH_DURING_RESET                                               -  60168 -  AWVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                     
// AXI_WVALID_HIGH_DURING_RESET                                                -  60169 -  WVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                       
// AXI_BVALID_HIGH_DURING_RESET                                                -  60170 -  BVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                        
// AXI_ARVALID_HIGH_DURING_RESET                                               -  60171 -  ARVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                          
// AXI_RVALID_HIGH_DURING_RESET                                                -  60172 -  RVALID asserted during the reset state (SPEC3(A3.1.2))                                                                                                                         
// AXI_RLAST_VIOLATION                                                         -  60173 -  RLAST signal should be asserted along with the final transfer of the read data burst (SPEC3(A3.4.1))                                                                                    
// AXI_EX_WRITE_AFTER_EX_READ_FAILURE                                          -  60174 -  It is recommended that an exclusive write access should not be performed after the corresponding exclusive read failure. (SPEC3(A7.2.2))                                
// AXI_TIMEOUT_WAITING_FOR_WRITE_DATA                                          -  60175 -  Timed-out waiting for a data phase in write data burst. SPEC3(A2.3)                                                           
// AXI_TIMEOUT_WAITING_FOR_WRITE_RESPONSE                                      -  60176 -  Timed-out waiting for a write response. SPEC3(A2.4)                                                                      
// AXI_TIMEOUT_WAITING_FOR_READ_RESPONSE                                       -  60177 -  Timed-out waiting for a read response. SPEC3(A2.6)                                                                            
// AXI_TIMEOUT_WAITING_FOR_WRITE_ADDR_AFTER_DATA                               -  60178 -  Timed-out waiting for a write address phase to be coming after data SPEC3(A2.2)                                       
// AXI_DEC_ERR_RESP_FOR_READ                                                   -  60179 -  No slave at the address for this read transfer (signaled by ~AXI_DECERR~)                                                                     
// AXI_DEC_ERR_RESP_FOR_WRITE                                                  -  60180 -  No slave at the address for this write transfer (signaled by ~AXI_DECERR~)                                                                     
// AXI_SLV_ERR_RESP_FOR_READ                                                   -  60181 -  Slave has detected an error for this read transfer (signaled by ~AXI_SLVERR~)                                                                  
// AXI_SLV_ERR_RESP_FOR_WRITE                                                  -  60182 -  Slave has detected an error for this write transfer (signaled by ~AXI_SLVERR~)                                                                   
// AXI_MINIMUM_SLAVE_ADDRESS_SPACE_VIOLATION                                   -  60183 -  The minimum address space occupied by a single slave device is 4 kilobytes (SPEC3(A10.3.2))                                       
// AXI_ADDRESS_WIDTH_EXCEEDS_64                                                -  60184 -  AXI supports up to 64-bit addressing (SPEC3(A10.3.1))                                                                                                                  
// AXI_READ_BURST_MAXIMUM_LENGTH_VIOLATION                                     -  60185 -  16 read data beats were seen without RLAST (SPEC3(A3.4.1))                                                                                                   
// AXI_WRITE_BURST_MAXIMUM_LENGTH_VIOLATION                                    -  60186 -  16 write data beats were seen without WLAST (see AMBA AXI and ACE Protocol Specification IHI0022D section A3.4.1 )                                     
// AXI_WRITE_STROBES_LENGTH_VIOLATION                                          -  60187 -  The size of the write_strobes array in a write transfer should match the value given by AWLEN                                                                                               
// AXI_EX_RD_WHEN_EX_NOT_ENABLED                                               -  60188 -  An exclusive read should not be issued when exclusive transactions are not enabled                                                                                                                   
// AXI_EX_WR_WHEN_EX_NOT_ENABLED                                               -  60189 -  An exclusive write should not be issued when exclusive transactions are not enabled                                                                                                     
// AXI_WRITE_TRANSFER_EXCEEDS_ADDRESS_SPACE                                    -  60190 -  This write transfer runs off the edge of the address space defined by AXI_ADDRESS_WIDTH (SPEC3(A10.3.1))                                                                           
// AXI_READ_TRANSFER_EXCEEDS_ADDRESS_SPACE                                     -  60191 -  This read transfer runs off the edge of the address space defined by AXI_ADDRESS_WIDTH (SPEC3(A10.3.1))                                                                                 
// AXI_EXCL_RD_WHILE_EXCL_WR_IN_PROGRESS_SAME_ID                               -  60192 -  Master starts an exclusive read burst while exclusive write burst with same ID tag is in progress (SPEC3(A7.2.4))                                                                 
// AXI_EXCL_WR_WHILE_EXCL_RD_IN_PROGRESS_SAME_ID                               -  60193 -  Master starts an exclusive write burst while exclusive read burst with same ID tag is in progress (SPEC3(A7.2.4))                                                                
// AXI_ILLEGAL_LENGTH_READ_BURST                                               -  60194 -  Read address phase burst_length has an illegal value (SPEC3(A3.4.1))                                                                                                                      
// AXI_ILLEGAL_LENGTH_WRITE_BURST                                              -  60195 -  Write address phase burst_length has an illegal value (SPEC3(A3.4.1))                                                                                                                        
// AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID                                      -  60196 -  Once ARVALID has been asserted, ARREADY> should be asserted within config_max_latency_ARVALID_assertion_to_ARREADY clock periods                                                     
// AXI_BREADY_NOT_ASSERTED_AFTER_BVALID                                        -  60197 -  Once BVALID has been asserted, BREADY> should be asserted within config_max_latency_BVALID_assertion_to_BREADY clock periods                                                             
// AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID                                      -  60198 -  Once AWVALID has been asserted, AWREADY> should be asserted within config_max_latency_AWVALID_assertion_to_AWREADY clock periods                                                              
// AXI_RREADY_NOT_ASSERTED_AFTER_RVALID                                        -  60199 -  Once RVALID has been asserted, RREADY> should be asserted within config_max_latency_RVALID_assertion_to_RREADY clock periods                                                                
// AXI_WREADY_NOT_ASSERTED_AFTER_WVALID                                        -  60200 -  Once WVALID has been asserted, WREADY> should be asserted within config_max_latency_WVALID_assertion_to_WREADY clock periods                                                           
// AXI_DEC_ERR_ILLEGAL_FOR_MAPPED_SLAVE_ADDR                                   -  60201 -  Slave receives a burst to a mapped address but responds with DECERR (signalled by AXI_DECERR) (SPEC3(A3.4.4))                                                                           
// AXI_PARAM_READ_REORDERING_DEPTH_EQUALS_ZERO                                 -  60202 -  The user-supplied config_read_data_reordering_depth should be greater than zero (SPEC3(A5.3.1))                                                                                        
// AXI_PARAM_READ_REORDERING_DEPTH_EXCEEDS_MAX_ID                              -  60203 -  The user-supplied config_read_data_reordering_depth exceeds the maximum possible value, as defined by the AXI_ID_WIDTH parameter (SPEC3(A5.3.1))                              
// AXI_READ_REORDERING_VIOLATION                                               -  60204 -  The arrival of a read response has exceeded the read reordering depth (SPEC3(A5.3.1))                             
// AXI_READ_ISSUING_CAPABILITY_VIOLATION                                       -  60205 -  Number of outstanding Read transactions exceeded maximum Read issuing capability 
// AXI_WRITE_ISSUING_CAPABILITY_VIOLATION                                      -  60206 -  Number of outstanding Write transactions exceeded maximum Write issuing capability
// AXI_COMBINED_ISSUING_CAPABILITY_VIOLATION                                   -  60207 -  Number of outstanding Read and Write transactions exceeded maximum combined issuing capability 
// AXI_READ_ACCEPTANCE_CAPABILITY_VIOLATION                                    -  60208 -  Number of outstanding Read transactions exceeded maximum Read acceptance capability 
// AXI_WRITE_ACCEPTANCE_CAPABILITY_VIOLATION                                   -  60209 -  Number of outstanding Write transactions exceeded maximum Write acceptance capability 
// AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION                                -  60210 -  Number of outstanding Read and Write transactions exceeded maximum combined acceptance capability 
typedef enum bit [7:0]
{
    AXI_ARESETn_SIGNAL_Z                                                        = 8'h00,
    AXI_ARESETn_SIGNAL_X                                                        = 8'h01,
    AXI_ACLK_SIGNAL_Z                                                           = 8'h02,
    AXI_ACLK_SIGNAL_X                                                           = 8'h03,
    AXI_ADDR_FOR_READ_BURST_ACROSS_4K_BOUNDARY                                  = 8'h04,
    AXI_ADDR_FOR_WRITE_BURST_ACROSS_4K_BOUNDARY                                 = 8'h05,
    AXI_ARADDR_CHANGED_BEFORE_ARREADY                                           = 8'h06,
    AXI_ARADDR_UNKN                                                             = 8'h07,
    AXI_ARBURST_CHANGED_BEFORE_ARREADY                                          = 8'h08,
    AXI_ARBURST_UNKN                                                            = 8'h09,
    AXI_ARCACHE_CHANGED_BEFORE_ARREADY                                          = 8'h0a,
    AXI_ARCACHE_UNKN                                                            = 8'h0b,
    AXI_ARID_CHANGED_BEFORE_ARREADY                                             = 8'h0c,
    AXI_ARID_UNKN                                                               = 8'h0d,
    AXI_ARLEN_CHANGED_BEFORE_ARREADY                                            = 8'h0e,
    AXI_ARLEN_UNKN                                                              = 8'h0f,
    AXI_ARLOCK_CHANGED_BEFORE_ARREADY                                           = 8'h10,
    AXI_ARLOCK_UNKN                                                             = 8'h11,
    AXI_ARPROT_CHANGED_BEFORE_ARREADY                                           = 8'h12,
    AXI_ARPROT_UNKN                                                             = 8'h13,
    AXI_ARREADY_UNKN                                                            = 8'h14,
    AXI_ARSIZE_CHANGED_BEFORE_ARREADY                                           = 8'h15,
    AXI_ARSIZE_UNKN                                                             = 8'h16,
    AXI_ARUSER_CHANGED_BEFORE_ARREADY                                           = 8'h17,
    AXI_ARUSER_UNKN                                                             = 8'h18,
    AXI_ARVALID_DEASSERTED_BEFORE_ARREADY                                       = 8'h19,
    AXI_ARVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                 = 8'h1a,
    AXI_ARVALID_UNKN                                                            = 8'h1b,
    AXI_AWADDR_CHANGED_BEFORE_AWREADY                                           = 8'h1c,
    AXI_AWADDR_UNKN                                                             = 8'h1d,
    AXI_AWBURST_CHANGED_BEFORE_AWREADY                                          = 8'h1e,
    AXI_AWBURST_UNKN                                                            = 8'h1f,
    AXI_AWCACHE_CHANGED_BEFORE_AWREADY                                          = 8'h20,
    AXI_AWCACHE_UNKN                                                            = 8'h21,
    AXI_AWID_CHANGED_BEFORE_AWREADY                                             = 8'h22,
    AXI_AWID_UNKN                                                               = 8'h23,
    AXI_AWLEN_CHANGED_BEFORE_AWREADY                                            = 8'h24,
    AXI_AWLEN_UNKN                                                              = 8'h25,
    AXI_AWLOCK_CHANGED_BEFORE_AWREADY                                           = 8'h26,
    AXI_AWLOCK_UNKN                                                             = 8'h27,
    AXI_AWPROT_CHANGED_BEFORE_AWREADY                                           = 8'h28,
    AXI_AWPROT_UNKN                                                             = 8'h29,
    AXI_AWREADY_UNKN                                                            = 8'h2a,
    AXI_AWSIZE_CHANGED_BEFORE_AWREADY                                           = 8'h2b,
    AXI_AWSIZE_UNKN                                                             = 8'h2c,
    AXI_AWUSER_CHANGED_BEFORE_AWREADY                                           = 8'h2d,
    AXI_AWUSER_UNKN                                                             = 8'h2e,
    AXI_AWVALID_DEASSERTED_BEFORE_AWREADY                                       = 8'h2f,
    AXI_AWVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                 = 8'h30,
    AXI_AWVALID_UNKN                                                            = 8'h31,
    AXI_BID_CHANGED_BEFORE_BREADY                                               = 8'h32,
    AXI_BID_UNKN                                                                = 8'h33,
    AXI_BREADY_UNKN                                                             = 8'h34,
    AXI_BRESP_CHANGED_BEFORE_BREADY                                             = 8'h35,
    AXI_BRESP_UNKN                                                              = 8'h36,
    AXI_BUSER_CHANGED_BEFORE_BREADY                                             = 8'h37,
    AXI_BUSER_UNKN                                                              = 8'h38,
    AXI_BVALID_DEASSERTED_BEFORE_BREADY                                         = 8'h39,
    AXI_BVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  = 8'h3a,
    AXI_BVALID_UNKN                                                             = 8'h3b,
    AXI_EXCLUSIVE_READ_ACCESS_MODIFIABLE                                        = 8'h3c,
    AXI_EXCLUSIVE_READ_BYTES_TRANSFER_EXCEEDS_128                               = 8'h3d,
    AXI_EXCLUSIVE_WRITE_BYTES_TRANSFER_EXCEEDS_128                              = 8'h3e,
    AXI_EXCLUSIVE_READ_BYTES_TRANSFER_NOT_POWER_OF_2                            = 8'h3f,
    AXI_EXCLUSIVE_WRITE_BYTES_TRANSFER_NOT_POWER_OF_2                           = 8'h40,
    AXI_EXCLUSIVE_WR_ADDRESS_NOT_SAME_AS_RD                                     = 8'h41,
    AXI_EXCLUSIVE_WR_BURST_NOT_SAME_AS_RD                                       = 8'h42,
    AXI_EXCLUSIVE_WR_CACHE_NOT_SAME_AS_RD                                       = 8'h43,
    AXI_EXCLUSIVE_WRITE_ACCESS_MODIFIABLE                                       = 8'h44,
    AXI_EXCLUSIVE_WR_LENGTH_NOT_SAME_AS_RD                                      = 8'h45,
    AXI_EXCLUSIVE_WR_PROT_NOT_SAME_AS_RD                                        = 8'h46,
    AXI_EXCLUSIVE_WR_SIZE_NOT_SAME_AS_RD                                        = 8'h47,
    AXI_EXOKAY_RESPONSE_NORMAL_READ                                             = 8'h48,
    AXI_EXOKAY_RESPONSE_NORMAL_WRITE                                            = 8'h49,
    AXI_EX_RD_RESP_MISMATCHED_WITH_EXPECTED_RESP                                = 8'h4a,
    AXI_EX_WR_RESP_MISMATCHED_WITH_EXPECTED_RESP                                = 8'h4b,
    AXI_EX_RD_EXOKAY_RESP_SLAVE_WITHOUT_EXCLUSIVE_ACCESS                        = 8'h4c,
    AXI_EX_WRITE_BEFORE_EX_READ_RESPONSE                                        = 8'h4d,
    AXI_EX_WRITE_EXOKAY_RESP_SLAVE_WITHOUT_EXCLUSIVE_ACCESS                     = 8'h4e,
    AXI_ILLEGAL_LENGTH_WRAPPING_READ_BURST                                      = 8'h4f,
    AXI_ILLEGAL_LENGTH_WRAPPING_WRITE_BURST                                     = 8'h50,
    AXI_ILLEGAL_RESPONSE_EXCLUSIVE_READ                                         = 8'h51,
    AXI_ILLEGAL_RESPONSE_EXCLUSIVE_WRITE                                        = 8'h52,
    AXI_PARAM_READ_DATA_BUS_WIDTH                                               = 8'h53,
    AXI_PARAM_WRITE_DATA_BUS_WIDTH                                              = 8'h54,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_12                                    = 8'h55,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_13                                    = 8'h56,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_4                                     = 8'h57,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_5                                     = 8'h58,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_8                                     = 8'h59,
    AXI_READ_ALLOCATE_WHEN_NON_MODIFIABLE_9                                     = 8'h5a,
    AXI_READ_BURST_LENGTH_VIOLATION                                             = 8'h5b,
    AXI_READ_BURST_SIZE_VIOLATION                                               = 8'h5c,
    AXI_READ_DATA_BEFORE_ADDRESS                                                = 8'h5d,
    AXI_READ_DATA_CHANGED_BEFORE_RREADY                                         = 8'h5e,
    AXI_READ_DATA_UNKN                                                          = 8'h5f,
    AXI_RESERVED_ARLOCK_ENCODING                                                = 8'h60,
    AXI_READ_RESP_CHANGED_BEFORE_RREADY                                         = 8'h61,
    AXI_RESERVED_ARBURST_ENCODING                                               = 8'h62,
    AXI_RESERVED_AWBURST_ENCODING                                               = 8'h63,
    AXI_RID_CHANGED_BEFORE_RREADY                                               = 8'h64,
    AXI_RID_UNKN                                                                = 8'h65,
    AXI_RLAST_CHANGED_BEFORE_RREADY                                             = 8'h66,
    AXI_RLAST_UNKN                                                              = 8'h67,
    AXI_RREADY_UNKN                                                             = 8'h68,
    AXI_RRESP_UNKN                                                              = 8'h69,
    AXI_RUSER_CHANGED_BEFORE_RREADY                                             = 8'h6a,
    AXI_RUSER_UNKN                                                              = 8'h6b,
    AXI_RVALID_DEASSERTED_BEFORE_RREADY                                         = 8'h6c,
    AXI_RVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  = 8'h6d,
    AXI_RVALID_UNKN                                                             = 8'h6e,
    AXI_UNALIGNED_ADDRESS_FOR_EXCLUSIVE_READ                                    = 8'h6f,
    AXI_UNALIGNED_ADDRESS_FOR_EXCLUSIVE_WRITE                                   = 8'h70,
    AXI_UNALIGNED_ADDR_FOR_WRAPPING_READ_BURST                                  = 8'h71,
    AXI_UNALIGNED_ADDR_FOR_WRAPPING_WRITE_BURST                                 = 8'h72,
    AXI_WDATA_CHANGED_BEFORE_WREADY_ON_INVALID_LANE                             = 8'h73,
    AXI_WDATA_CHANGED_BEFORE_WREADY_ON_VALID_LANE                               = 8'h74,
    AXI_WLAST_CHANGED_BEFORE_WREADY                                             = 8'h75,
    AXI_WID_CHANGED_BEFORE_WREADY                                               = 8'h76,
    AXI_WLAST_UNKN                                                              = 8'h77,
    AXI_WID_UNKN                                                                = 8'h78,
    AXI_WREADY_UNKN                                                             = 8'h79,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_12                                   = 8'h7a,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_13                                   = 8'h7b,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_4                                    = 8'h7c,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_5                                    = 8'h7d,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_8                                    = 8'h7e,
    AXI_WRITE_ALLOCATE_WHEN_NON_MODIFIABLE_9                                    = 8'h7f,
    AXI_WRITE_BURST_SIZE_VIOLATION                                              = 8'h80,
    AXI_WRITE_DATA_BEFORE_ADDRESS                                               = 8'h81,
    AXI_WRITE_DATA_UNKN_ON_INVALID_LANE                                         = 8'h82,
    AXI_WRITE_DATA_UNKN_ON_VALID_LANE                                           = 8'h83,
    AXI_RESERVED_AWLOCK_ENCODING                                                = 8'h84,
    AXI_WRITE_STROBE_ON_INVALID_BYTE_LANES                                      = 8'h85,
    AXI_WSTRB_CHANGED_BEFORE_WREADY                                             = 8'h86,
    AXI_WSTRB_UNKN                                                              = 8'h87,
    AXI_WUSER_CHANGED_BEFORE_WREADY                                             = 8'h88,
    AXI_WUSER_UNKN                                                              = 8'h89,
    AXI_WVALID_DEASSERTED_BEFORE_WREADY                                         = 8'h8a,
    AXI_WVALID_HIGH_ON_FIRST_CLOCK_AFTER_RESET                                  = 8'h8b,
    AXI_WVALID_UNKN                                                             = 8'h8c,
    AXI_ADDR_ACROSS_4K_WITHIN_LOCKED_WRITE_TRANSACTION                          = 8'h8d,
    AXI_ADDR_ACROSS_4K_WITHIN_LOCKED_READ_TRANSACTION                           = 8'h8e,
    AXI_AWID_CHANGED_WITHIN_LOCKED_TRANSACTION                                  = 8'h8f,
    AXI_ARID_CHANGED_WITHIN_LOCKED_TRANSACTION                                  = 8'h90,
    AXI_AWPROT_CHANGED_WITHIN_LOCKED_TRANSACTION                                = 8'h91,
    AXI_ARPROT_CHANGED_WITHIN_LOCKED_TRANSACTION                                = 8'h92,
    AXI_AWCACHE_CHANGED_WITHIN_LOCKED_TRANSACTION                               = 8'h93,
    AXI_ARCACHE_CHANGED_WITHIN_LOCKED_TRANSACTION                               = 8'h94,
    AXI_NUMBER_OF_LOCKED_SEQUENCES_EXCEEDS_2                                    = 8'h95,
    AXI_LOCKED_WRITE_BEFORE_COMPLETION_OF_PREVIOUS_WRITE_TRANSACTIONS           = 8'h96,
    AXI_LOCKED_WRITE_BEFORE_COMPLETION_OF_PREVIOUS_READ_TRANSACTIONS            = 8'h97,
    AXI_LOCKED_READ_BEFORE_COMPLETION_OF_PREVIOUS_WRITE_TRANSACTIONS            = 8'h98,
    AXI_LOCKED_READ_BEFORE_COMPLETION_OF_PREVIOUS_READ_TRANSACTIONS             = 8'h99,
    AXI_NEW_BURST_BEFORE_COMPLETION_OF_UNLOCK_TRANSACTION                       = 8'h9a,
    AXI_UNLOCKED_WRITE_WHILE_OUTSTANDING_LOCKED_WRITES                          = 8'h9b,
    AXI_UNLOCKED_WRITE_WHILE_OUTSTANDING_LOCKED_READS                           = 8'h9c,
    AXI_UNLOCKED_READ_WHILE_OUTSTANDING_LOCKED_WRITES                           = 8'h9d,
    AXI_UNLOCKED_READ_WHILE_OUTSTANDING_LOCKED_READS                            = 8'h9e,
    AXI_UNLOCKING_TRANSACTION_WITH_AN_EXCLUSIVE_ACCESS                          = 8'h9f,
    AXI_FIRST_DATA_ITEM_OF_TRANSACTION_WRITE_ORDER_VIOLATION                    = 8'ha0,
    AXI_AWLEN_MISMATCHED_WITH_COMPLETED_WRITE_DATA_BURST                        = 8'ha1,
    AXI_WRITE_LENGTH_MISMATCHED_ACTUAL_LENGTH_OF_WRITE_DATA_BURST_EXCEEDS_AWLEN = 8'ha2,
    AXI_AWLEN_MISMATCHED_ACTUAL_LENGTH_OF_WRITE_DATA_BURST_EXCEEDS_AWLEN        = 8'ha3,
    AXI_WLAST_ASSERTED_DURING_DATA_PHASE_OTHER_THAN_LAST                        = 8'ha4,
    AXI_WRITE_INTERLEAVE_DEPTH_VIOLATION                                        = 8'ha5,
    AXI_WRITE_RESPONSE_WITHOUT_ADDR                                             = 8'ha6,
    AXI_WRITE_RESPONSE_WITHOUT_DATA                                             = 8'ha7,
    AXI_AWVALID_HIGH_DURING_RESET                                               = 8'ha8,
    AXI_WVALID_HIGH_DURING_RESET                                                = 8'ha9,
    AXI_BVALID_HIGH_DURING_RESET                                                = 8'haa,
    AXI_ARVALID_HIGH_DURING_RESET                                               = 8'hab,
    AXI_RVALID_HIGH_DURING_RESET                                                = 8'hac,
    AXI_RLAST_VIOLATION                                                         = 8'had,
    AXI_EX_WRITE_AFTER_EX_READ_FAILURE                                          = 8'hae,
    AXI_TIMEOUT_WAITING_FOR_WRITE_DATA                                          = 8'haf,
    AXI_TIMEOUT_WAITING_FOR_WRITE_RESPONSE                                      = 8'hb0,
    AXI_TIMEOUT_WAITING_FOR_READ_RESPONSE                                       = 8'hb1,
    AXI_TIMEOUT_WAITING_FOR_WRITE_ADDR_AFTER_DATA                               = 8'hb2,
    AXI_DEC_ERR_RESP_FOR_READ                                                   = 8'hb3,
    AXI_DEC_ERR_RESP_FOR_WRITE                                                  = 8'hb4,
    AXI_SLV_ERR_RESP_FOR_READ                                                   = 8'hb5,
    AXI_SLV_ERR_RESP_FOR_WRITE                                                  = 8'hb6,
    AXI_MINIMUM_SLAVE_ADDRESS_SPACE_VIOLATION                                   = 8'hb7,
    AXI_ADDRESS_WIDTH_EXCEEDS_64                                                = 8'hb8,
    AXI_READ_BURST_MAXIMUM_LENGTH_VIOLATION                                     = 8'hb9,
    AXI_WRITE_BURST_MAXIMUM_LENGTH_VIOLATION                                    = 8'hba,
    AXI_WRITE_STROBES_LENGTH_VIOLATION                                          = 8'hbb,
    AXI_EX_RD_WHEN_EX_NOT_ENABLED                                               = 8'hbc,
    AXI_EX_WR_WHEN_EX_NOT_ENABLED                                               = 8'hbd,
    AXI_WRITE_TRANSFER_EXCEEDS_ADDRESS_SPACE                                    = 8'hbe,
    AXI_READ_TRANSFER_EXCEEDS_ADDRESS_SPACE                                     = 8'hbf,
    AXI_EXCL_RD_WHILE_EXCL_WR_IN_PROGRESS_SAME_ID                               = 8'hc0,
    AXI_EXCL_WR_WHILE_EXCL_RD_IN_PROGRESS_SAME_ID                               = 8'hc1,
    AXI_ILLEGAL_LENGTH_READ_BURST                                               = 8'hc2,
    AXI_ILLEGAL_LENGTH_WRITE_BURST                                              = 8'hc3,
    AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID                                      = 8'hc4,
    AXI_BREADY_NOT_ASSERTED_AFTER_BVALID                                        = 8'hc5,
    AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID                                      = 8'hc6,
    AXI_RREADY_NOT_ASSERTED_AFTER_RVALID                                        = 8'hc7,
    AXI_WREADY_NOT_ASSERTED_AFTER_WVALID                                        = 8'hc8,
    AXI_DEC_ERR_ILLEGAL_FOR_MAPPED_SLAVE_ADDR                                   = 8'hc9,
    AXI_PARAM_READ_REORDERING_DEPTH_EQUALS_ZERO                                 = 8'hca,
    AXI_PARAM_READ_REORDERING_DEPTH_EXCEEDS_MAX_ID                              = 8'hcb,
    AXI_READ_REORDERING_VIOLATION                                               = 8'hcc,
    AXI_READ_ISSUING_CAPABILITY_VIOLATION                                       = 8'hcd,
    AXI_WRITE_ISSUING_CAPABILITY_VIOLATION                                      = 8'hce,
    AXI_COMBINED_ISSUING_CAPABILITY_VIOLATION                                   = 8'hcf,
    AXI_READ_ACCEPTANCE_CAPABILITY_VIOLATION                                    = 8'hd0,
    AXI_WRITE_ACCEPTANCE_CAPABILITY_VIOLATION                                   = 8'hd1,
    AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION                                = 8'hd2
} axi_assertion_e;



//------------------------------------------------------------------------------
//
// Enum: axi_ready_e
//
//------------------------------------------------------------------------------
// 
//  Specifies wait if AXI_NOT_READY and specifies no wait if AXI_READY.
// 
typedef enum bit [0:0]
{
    AXI_NOT_READY = 1'h0,
    AXI_READY     = 1'h1
} axi_ready_e;



//------------------------------------------------------------------------------
//
// Enum: axi_wtrans_phase_e
//
//------------------------------------------------------------------------------
// 
//  An enumerated type used in the coverage collector class
//  <axi_functional_coverage> for encoding the address/data/response type for each
//  phase of a write transaction.
// 
//  As each phase of a write occurs, a field of the <axi_write_trans_record>
//  record is updated with the type (address/data/response) of the phase (this
//  information is used at the end of the transaction to classify the
//  <axi_functional_coverage::axi_wtrans_phase_order_e> phase-ordering type of the
//  transaction).
//  See the <axi_functional_coverage::put_wphase> task.
// 
//  A (ADDR) - The address phase of a write transaction.
//  D (DATA) - The data phase of a write transaction.
//  R (RESP) - The response phase of a write transaction.
// 
typedef enum bit [1:0]
{
    A = 2'h0,
    D = 2'h1,
    R = 2'h2
} axi_wtrans_phase_e;


//------------------------------------------------------------------------------
//
// Struct: axi_rw_txn_counts_s
//
//------------------------------------------------------------------------------

typedef struct packed
{
    int unsigned reads_no_resp;
    int unsigned reads_no_resp_for_id;
    int unsigned waddr_no_resp;
    int unsigned waddr_no_resp_for_id;
    int unsigned wdata_no_resp;
    int unsigned wdata_no_resp_for_id;
    int unsigned writes_no_resp;
    int unsigned writes_no_resp_for_id;
} axi_rw_txn_counts_s;



typedef bit [1023:0] axi_max_bits_t;

// enum: axi_config_e
//
// An enum which fields corresponding to each configuration parameter of the VIP
//    AXI_CONFIG_WRITE_CTRL_TO_DATA_MINTIME - 
//         
//         Sets the delay from start of address phase to start of data phase in a write 
//         transaction (in terms of ACLK).
//         
//         Default: 1 
//         
//         This configuration variable has been deprecated and is maintained 
//         for backward compatibility. However, you can use ~write_address_to_data_delay~ 
//         configuration variable to control the delay between a write address phase 
//         and a write data phase.
//         
//    AXI_CONFIG_ENABLE_ALL_ASSERTIONS - 
//         
//         Enables all protocol assertions. 
//         
//         Default: 1
//         
//    AXI_CONFIG_ENABLE_ASSERTION - 
//         
//         Enables individual protocol assertion.
//         This variable controls whether specific assertion within QVIP (of type <axi_assertion_e>) is enabled or disabled.
//         Individual assertion can be disabled as follows:-
//         //-----------------------------------------------------------------------
//         // < BFM interface>.set_config_enable_assertion_index1(<name of assertion>,1'b0);
//         //-----------------------------------------------------------------------
//         
//         For example, the assertion AXI_READ_DATA_UNKN is disabled as follows:
//         <bfm>.set_config_enable_assertion_index1(AXI_READ_DATA_UNKN, 1'b0); 
//         
//         Here bfm is the AXI interface instance name for which the assertion to be disabled. 
//         
//         Default: All assertions are enabled
//           
//         
//    AXI_CONFIG_SUPPORT_EXCLUSIVE_ACCESS - 
//         
//         Enables exclusive transactions support for slave.
//         If disabled, every exclusive read/write returns an OKAY response,
//         and exclusive write updates memory. 
//         
//         Default: 1  
//         
//    AXI_CONFIG_READ_DATA_REORDERING_DEPTH - 
//         
//         Sets the maximum number of different read transaction addresses for which read 
//         data(response) can be sent in any order from slave. 
//         
//         Default: 2 ** AXI_ID_WIDTH
//         
//    AXI_CONFIG_MAX_TRANSACTION_TIME_FACTOR - 
//          
//         Sets maximum timeout period (in terms of ACLK) for any complete read or write transaction, which
//         includes time period for all individual phases of transaction. 
//         
//         Default: 100000 clock cycles
//         
//    AXI_CONFIG_TIMEOUT_MAX_DATA_TRANSFER - 
//          
//         Sets maximum number of write data beats in a write data burst. 
//         
//         Default: 1024  
//         
//    AXI_CONFIG_BURST_TIMEOUT_FACTOR - 
//          
//         Sets maximum timeout period (in terms of ACLK) between individual phases of a transaction. 
//         
//         Default: 10000 clock cycles 
//         
//    AXI_CONFIG_MAX_LATENCY_AWVALID_ASSERTION_TO_AWREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of AWVALID to assertion of AWREADY.
//         An error message AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID is generated if AWREADY is not asserted
//         after assertion of AWVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MAX_LATENCY_ARVALID_ASSERTION_TO_ARREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of ARVALID to assertion of ARREADY.
//         An error message AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID is generated if ARREADY is not asserted
//         after assertion of ARVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MAX_LATENCY_RVALID_ASSERTION_TO_RREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of RVALID to assertion of RREADY.
//         An error message AXI_RREADY_NOT_ASSERTED_AFTER_RVALID is generated if RREADY is not asserted
//         after assertion of RVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MAX_LATENCY_BVALID_ASSERTION_TO_BREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of BVALID to assertion of BREADY.
//         An error message AXI_BREADY_NOT_ASSERTED_AFTER_BVALID is generated if BREADY is not asserted
//         after assertion of BVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MAX_LATENCY_WVALID_ASSERTION_TO_WREADY - 
//          
//         Sets maximum timeout period (in terms of ACLK) from assertion of WVALID to assertion of WREADY.
//         An error message AXI_WREADY_NOT_ASSERTED_AFTER_WVALID is generated if WREADY is not asserted
//         after assertion of WVALID within this period. 
//         
//         Default: 10000 clock cycles
//         
//    AXI_CONFIG_MASTER_ERROR_POSITION - 
//         
//         Sets type of master error.
//         
//    AXI_CONFIG_SETUP_TIME - 
//         
//         Sets number of simulation time units from the setup time to the active 
//         clock edge of ACLK. The setup time will always be less than the time period
//         of the clock. 
//         
//         Default: 0
//         
//    AXI_CONFIG_HOLD_TIME - 
//         
//         Sets number of simulation time units from the hold time to the active 
//         clock edge of ACLK. 
//         
//         Default: 0
//         
//    AXI_CONFIG_MAX_OUTSTANDING_WR -  Configures maximum possible outstanding Write transactions
//    AXI_CONFIG_MAX_OUTSTANDING_RD -  Configures maximum possible outstanding Read transactions
//    AXI_CONFIG_MAX_OUTSTANDING_RW -  Configures maximum possible outstanding Combined (Read and Write) transactions
//    AXI_CONFIG_IS_ISSUING -  Enables Master component to use "config_max_outstanding_wr/config_max_outstanding_rd/config_max_outstanding_rw" variables for transaction issuing capability when set to true

typedef enum bit [7:0]
{
    AXI_CONFIG_WRITE_CTRL_TO_DATA_MINTIME    = 8'd0,
    AXI_CONFIG_MASTER_WRITE_DELAY            = 8'd1,
    AXI_CONFIG_ENABLE_ALL_ASSERTIONS         = 8'd2,
    AXI_CONFIG_ENABLE_ASSERTION              = 8'd3,
    AXI_CONFIG_SLAVE_START_ADDR              = 8'd4,
    AXI_CONFIG_SLAVE_END_ADDR                = 8'd5,
    AXI_CONFIG_SUPPORT_EXCLUSIVE_ACCESS      = 8'd6,
    AXI_CONFIG_READ_DATA_REORDERING_DEPTH    = 8'd7,
    AXI_CONFIG_MAX_TRANSACTION_TIME_FACTOR   = 8'd8,
    AXI_CONFIG_TIMEOUT_MAX_DATA_TRANSFER     = 8'd9,
    AXI_CONFIG_BURST_TIMEOUT_FACTOR          = 8'd10,
    AXI_CONFIG_MAX_LATENCY_AWVALID_ASSERTION_TO_AWREADY = 8'd11,
    AXI_CONFIG_MAX_LATENCY_ARVALID_ASSERTION_TO_ARREADY = 8'd12,
    AXI_CONFIG_MAX_LATENCY_RVALID_ASSERTION_TO_RREADY = 8'd13,
    AXI_CONFIG_MAX_LATENCY_BVALID_ASSERTION_TO_BREADY = 8'd14,
    AXI_CONFIG_MAX_LATENCY_WVALID_ASSERTION_TO_WREADY = 8'd15,
    AXI_CONFIG_MASTER_ERROR_POSITION         = 8'd16,
    AXI_CONFIG_SETUP_TIME                    = 8'd17,
    AXI_CONFIG_HOLD_TIME                     = 8'd18,
    AXI_CONFIG_MAX_OUTSTANDING_WR            = 8'd19,
    AXI_CONFIG_MAX_OUTSTANDING_RD            = 8'd20,
    AXI_CONFIG_MAX_OUTSTANDING_RW            = 8'd21,
    AXI_CONFIG_IS_ISSUING                    = 8'd22
} axi_config_e;

// enum: axi_vhd_if_e
//
// For VHDL use only
typedef enum int
{
    AXI_VHD_SET_CONFIG                         = 32'd0,
    AXI_VHD_GET_CONFIG                         = 32'd1,
    AXI_VHD_CREATE_WRITE_TRANSACTION           = 32'd2,
    AXI_VHD_CREATE_READ_TRANSACTION            = 32'd3,
    AXI_VHD_SET_ADDR                           = 32'd4,
    AXI_VHD_GET_ADDR                           = 32'd5,
    AXI_VHD_SET_SIZE                           = 32'd6,
    AXI_VHD_GET_SIZE                           = 32'd7,
    AXI_VHD_SET_BURST                          = 32'd8,
    AXI_VHD_GET_BURST                          = 32'd9,
    AXI_VHD_SET_LOCK                           = 32'd10,
    AXI_VHD_GET_LOCK                           = 32'd11,
    AXI_VHD_SET_CACHE                          = 32'd12,
    AXI_VHD_GET_CACHE                          = 32'd13,
    AXI_VHD_SET_PROT                           = 32'd14,
    AXI_VHD_GET_PROT                           = 32'd15,
    AXI_VHD_SET_ID                             = 32'd16,
    AXI_VHD_GET_ID                             = 32'd17,
    AXI_VHD_SET_BURST_LENGTH                   = 32'd18,
    AXI_VHD_GET_BURST_LENGTH                   = 32'd19,
    AXI_VHD_SET_DATA_WORDS                     = 32'd20,
    AXI_VHD_GET_DATA_WORDS                     = 32'd21,
    AXI_VHD_SET_WRITE_STROBES                  = 32'd22,
    AXI_VHD_GET_WRITE_STROBES                  = 32'd23,
    AXI_VHD_SET_RESP                           = 32'd24,
    AXI_VHD_GET_RESP                           = 32'd25,
    AXI_VHD_SET_ADDR_USER                      = 32'd26,
    AXI_VHD_GET_ADDR_USER                      = 32'd27,
    AXI_VHD_SET_READ_OR_WRITE                  = 32'd28,
    AXI_VHD_GET_READ_OR_WRITE                  = 32'd29,
    AXI_VHD_SET_ADDRESS_VALID_DELAY            = 32'd30,
    AXI_VHD_GET_ADDRESS_VALID_DELAY            = 32'd31,
    AXI_VHD_SET_DATA_VALID_DELAY               = 32'd32,
    AXI_VHD_GET_DATA_VALID_DELAY               = 32'd33,
    AXI_VHD_SET_WRITE_RESPONSE_VALID_DELAY     = 32'd34,
    AXI_VHD_GET_WRITE_RESPONSE_VALID_DELAY     = 32'd35,
    AXI_VHD_SET_ADDRESS_READY_DELAY            = 32'd36,
    AXI_VHD_GET_ADDRESS_READY_DELAY            = 32'd37,
    AXI_VHD_SET_DATA_READY_DELAY               = 32'd38,
    AXI_VHD_GET_DATA_READY_DELAY               = 32'd39,
    AXI_VHD_SET_WRITE_RESPONSE_READY_DELAY     = 32'd40,
    AXI_VHD_GET_WRITE_RESPONSE_READY_DELAY     = 32'd41,
    AXI_VHD_SET_GEN_WRITE_STROBES              = 32'd42,
    AXI_VHD_GET_GEN_WRITE_STROBES              = 32'd43,
    AXI_VHD_SET_OPERATION_MODE                 = 32'd44,
    AXI_VHD_GET_OPERATION_MODE                 = 32'd45,
    AXI_VHD_SET_DELAY_MODE                     = 32'd46,
    AXI_VHD_GET_DELAY_MODE                     = 32'd47,
    AXI_VHD_SET_WRITE_DATA_MODE                = 32'd48,
    AXI_VHD_GET_WRITE_DATA_MODE                = 32'd49,
    AXI_VHD_SET_DATA_BEAT_DONE                 = 32'd50,
    AXI_VHD_GET_DATA_BEAT_DONE                 = 32'd51,
    AXI_VHD_SET_TRANSACTION_DONE               = 32'd52,
    AXI_VHD_GET_TRANSACTION_DONE               = 32'd53,
    AXI_VHD_EXECUTE_TRANSACTION                = 32'd54,
    AXI_VHD_GET_RW_TRANSACTION                 = 32'd55,
    AXI_VHD_EXECUTE_READ_DATA_BURST            = 32'd56,
    AXI_VHD_GET_READ_DATA_BURST                = 32'd57,
    AXI_VHD_EXECUTE_WRITE_DATA_BURST           = 32'd58,
    AXI_VHD_GET_WRITE_DATA_BURST               = 32'd59,
    AXI_VHD_EXECUTE_READ_ADDR_PHASE            = 32'd60,
    AXI_VHD_GET_READ_ADDR_PHASE                = 32'd61,
    AXI_VHD_EXECUTE_READ_DATA_PHASE            = 32'd62,
    AXI_VHD_GET_READ_DATA_PHASE                = 32'd63,
    AXI_VHD_EXECUTE_WRITE_ADDR_PHASE           = 32'd64,
    AXI_VHD_GET_WRITE_ADDR_PHASE               = 32'd65,
    AXI_VHD_EXECUTE_WRITE_DATA_PHASE           = 32'd66,
    AXI_VHD_GET_WRITE_DATA_PHASE               = 32'd67,
    AXI_VHD_EXECUTE_WRITE_RESPONSE_PHASE       = 32'd68,
    AXI_VHD_GET_WRITE_RESPONSE_PHASE           = 32'd69,
    AXI_VHD_CREATE_MONITOR_TRANSACTION         = 32'd70,
    AXI_VHD_CREATE_SLAVE_TRANSACTION           = 32'd71,
    AXI_VHD_PUSH_TRANSACTION_ID                = 32'd72,
    AXI_VHD_POP_TRANSACTION_ID                 = 32'd73,
    AXI_VHD_GET_WRITE_ADDR_DATA                = 32'd74,
    AXI_VHD_GET_READ_ADDR                      = 32'd75,
    AXI_VHD_SET_READ_DATA                      = 32'd76,
    AXI_VHD_PRINT                              = 32'd77,
    AXI_VHD_DESTRUCT_TRANSACTION               = 32'd78,
    AXI_VHD_WAIT_ON                            = 32'd79
} axi_vhd_if_e;


typedef enum bit [7:0]
{
    AXI_CLOCK_POSEDGE = 8'd0,
    AXI_CLOCK_NEGEDGE = 8'd1,
    AXI_CLOCK_ANYEDGE = 8'd2,
    AXI_CLOCK_0_TO_1  = 8'd3,
    AXI_CLOCK_1_TO_0  = 8'd4,
    AXI_RESET_POSEDGE = 8'd5,
    AXI_RESET_NEGEDGE = 8'd6,
    AXI_RESET_ANYEDGE = 8'd7,
    AXI_RESET_0_TO_1  = 8'd8,
    AXI_RESET_1_TO_0  = 8'd9
} axi_wait_e;

`ifndef MAX_AXI_ADDRESS_WIDTH
  `define MAX_AXI_ADDRESS_WIDTH 64
`endif

`ifndef MAX_AXI_RDATA_WIDTH
  `define MAX_AXI_RDATA_WIDTH 1024
`endif

`ifndef MAX_AXI_WDATA_WIDTH
  `define MAX_AXI_WDATA_WIDTH 1024
`endif

`ifndef MAX_AXI_ID_WIDTH
  `define MAX_AXI_ID_WIDTH 18
`endif

// enum: axi_operation_mode_e
//
typedef enum int
{
    AXI_TRANSACTION_NON_BLOCKING = 32'd0,
    AXI_TRANSACTION_BLOCKING     = 32'd1
} axi_operation_mode_e;

// enum: axi_delay_mode_e
//
typedef enum int
{
    AXI_VALID2READY = 32'd0,
    AXI_TRANS2READY = 32'd1
} axi_delay_mode_e;

// enum: axi_write_data_mode_e
//
typedef enum int
{
    AXI_DATA_AFTER_ADDRESS = 32'd0,
    AXI_DATA_WITH_ADDRESS  = 32'd1
} axi_write_data_mode_e;

// Global Transaction Class
class axi_transaction;
    // Protocol 
    bit [((`MAX_AXI_ADDRESS_WIDTH) - 1):0]  addr;
    axi_size_e size;
    axi_burst_e burst;
    axi_lock_e lock;
    axi_cache_e cache;
    axi_prot_e prot;
    bit [((`MAX_AXI_ID_WIDTH) - 1):0]  id;
    bit [3:0] burst_length;
    bit [((((`MAX_AXI_RDATA_WIDTH > `MAX_AXI_WDATA_WIDTH) ? `MAX_AXI_RDATA_WIDTH : `MAX_AXI_WDATA_WIDTH)) - 1):0] data_words [];
    bit [(((`MAX_AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [];
    axi_response_e resp[];
    bit [7:0] addr_user;
    axi_rw_e read_or_write;
    int address_valid_delay;
    int data_valid_delay[];
    int write_response_valid_delay;
    int address_ready_delay;
    int data_ready_delay[];
    int write_response_ready_delay;

    // Housekeeping
    bit gen_write_strobes = 1'b1;
    axi_operation_mode_e  operation_mode  = AXI_TRANSACTION_BLOCKING;
    axi_delay_mode_e      delay_mode      = AXI_VALID2READY;
    axi_write_data_mode_e write_data_mode = AXI_DATA_WITH_ADDRESS;
    bit data_beat_done[];
    bit transaction_done;

    // This varaible is for printing component name and should not be visible/documented
    string driver_name;

    function void set_addr( input bit [((`MAX_AXI_ADDRESS_WIDTH) - 1):0]  laddr );
      addr = laddr;
    endfunction

    function bit [((`MAX_AXI_ADDRESS_WIDTH) - 1):0]   get_addr();
      return addr;
    endfunction

    function void set_size( input axi_size_e lsize );
      size = lsize;
    endfunction

    function axi_size_e get_size();
      return size;
    endfunction

    function void set_burst( input axi_burst_e lburst );
      burst = lburst;
    endfunction

    function axi_burst_e get_burst();
      return burst;
    endfunction

    function void set_lock( input axi_lock_e llock );
      lock = llock;
    endfunction

    function axi_lock_e get_lock();
      return lock;
    endfunction

    function void set_cache( input axi_cache_e lcache );
      cache = lcache;
    endfunction

    function axi_cache_e get_cache();
      return cache;
    endfunction

    function void set_prot( input axi_prot_e lprot );
      prot = lprot;
    endfunction

    function axi_prot_e get_prot();
      return prot;
    endfunction

    function void set_id( input bit [((`MAX_AXI_ID_WIDTH) - 1):0]  lid );
      id = lid;
    endfunction

    function bit [((`MAX_AXI_ID_WIDTH) - 1):0]   get_id();
      return id;
    endfunction

    function void set_burst_length( input bit [3:0] lburst_length );
      burst_length = lburst_length;
      data_words           = new[(lburst_length + 1)];
      write_strobes        = new[(lburst_length + 1)];
      resp                 = new[(lburst_length + 1)];
      data_valid_delay     = new[(lburst_length + 1)];
      data_ready_delay     = new[(lburst_length + 1)];
      data_beat_done       = new[(lburst_length + 1)];
    endfunction

    function bit [3:0]  get_burst_length();
      return burst_length;
    endfunction

    function void set_data_words( input bit [((((`MAX_AXI_RDATA_WIDTH > `MAX_AXI_WDATA_WIDTH) ? `MAX_AXI_RDATA_WIDTH : `MAX_AXI_WDATA_WIDTH)) - 1):0] ldata_words, input int index = 0 );
      data_words[index] = ldata_words;
    endfunction

    function bit [((((`MAX_AXI_RDATA_WIDTH > `MAX_AXI_WDATA_WIDTH) ? `MAX_AXI_RDATA_WIDTH : `MAX_AXI_WDATA_WIDTH)) - 1):0]  get_data_words( input int index = 0 );
      return data_words[index];
    endfunction

    function void set_write_strobes( input bit [(((`MAX_AXI_WDATA_WIDTH / 8)) - 1):0] lwrite_strobes, input int index = 0 );
      write_strobes[index] = lwrite_strobes;
    endfunction

    function bit [(((`MAX_AXI_WDATA_WIDTH / 8)) - 1):0]  get_write_strobes( input int index = 0 );
      return write_strobes[index];
    endfunction

    function void set_resp( input axi_response_e lresp, input int index = 0 );
      resp[index] = lresp;
    endfunction

    function axi_response_e get_resp( input int index = 0 );
      return resp[index];
    endfunction

    function void set_addr_user( input bit [7:0] laddr_user );
      addr_user = laddr_user;
    endfunction

    function bit [7:0]  get_addr_user();
      return addr_user;
    endfunction

    function void set_read_or_write( input axi_rw_e lread_or_write );
      read_or_write = lread_or_write;
    endfunction

    function axi_rw_e get_read_or_write();
      return read_or_write;
    endfunction

    function void set_address_valid_delay( input int laddress_valid_delay );
      address_valid_delay = laddress_valid_delay;
    endfunction

    function int get_address_valid_delay();
      return address_valid_delay;
    endfunction

    function void set_data_valid_delay( input int ldata_valid_delay, input int index = 0 );
      data_valid_delay[index] = ldata_valid_delay;
    endfunction

    function int get_data_valid_delay( input int index = 0 );
      return data_valid_delay[index];
    endfunction

    function void set_write_response_valid_delay( input int lwrite_response_valid_delay );
      write_response_valid_delay = lwrite_response_valid_delay;
    endfunction

    function int get_write_response_valid_delay();
      return write_response_valid_delay;
    endfunction

    function void set_address_ready_delay( input int laddress_ready_delay );
      address_ready_delay = laddress_ready_delay;
    endfunction

    function int get_address_ready_delay();
      return address_ready_delay;
    endfunction

    function void set_data_ready_delay( input int ldata_ready_delay, input int index = 0 );
      data_ready_delay[index] = ldata_ready_delay;
    endfunction

    function int get_data_ready_delay( input int index = 0 );
      return data_ready_delay[index];
    endfunction

    function void set_write_response_ready_delay( input int lwrite_response_ready_delay );
      write_response_ready_delay = lwrite_response_ready_delay;
    endfunction

    function int get_write_response_ready_delay();
      return write_response_ready_delay;
    endfunction

    function void set_gen_write_strobes( input bit lgen_write_strobes);
      gen_write_strobes = lgen_write_strobes;
    endfunction

    function bit get_gen_write_strobes();
      return gen_write_strobes;
    endfunction

    function void set_operation_mode( input axi_operation_mode_e loperation_mode );
      operation_mode = loperation_mode;
    endfunction

    function axi_operation_mode_e get_operation_mode();
      return operation_mode;
    endfunction

    function void set_delay_mode( input axi_delay_mode_e ldelay_mode );
      delay_mode = ldelay_mode;
    endfunction

    function axi_delay_mode_e get_delay_mode();
      return delay_mode;
    endfunction

    function void set_write_data_mode( input axi_write_data_mode_e lwrite_data_mode );
      write_data_mode = lwrite_data_mode;
    endfunction

    function axi_write_data_mode_e get_write_data_mode();
      return write_data_mode;
    endfunction

    function void set_data_beat_done( input int ldata_beat_done, input int index = 0 );
      data_beat_done[index] = ldata_beat_done;
    endfunction

    function int get_data_beat_done( input int index = 0 );
      return data_beat_done[index];
    endfunction

    function void set_transaction_done( input int ltransaction_done );
      transaction_done = ltransaction_done;
    endfunction

    function int get_transaction_done();
      return transaction_done;
    endfunction

    // Function: do_print
    //
    // Prints axi_transaction transaction attributes
    function void print (bit print_delays = 1'b0);
      $display("------------------------------------------------------------------------");
      $display("%0t: %s axi_transaction", $time, driver_name);
      $display("------------------------------------------------------------------------");
      $display("addr : 'h%h", addr);
      $display("size : %s", size.name());
      $display("burst : %s", burst.name());
      $display("lock : %s", lock.name());
      $display("cache : %s", cache.name());
      $display("prot : %s", prot.name());
      $display("id : 'h%h", id);
      $display("burst_length : 'h%h", burst_length);
      foreach( data_words[i0_1] )
        $display("data_words[%0d] : 'h%h", i0_1, data_words[i0_1]);
      foreach( write_strobes[i0_1] )
        $display("write_strobes[%0d] : 'h%h", i0_1, write_strobes[i0_1]);
      foreach( resp[i0_1] )
        $display("resp[%0d] : %s", i0_1, resp[i0_1].name());
      $display("addr_user : 'h%h", addr_user);
      $display("read_or_write : %s", read_or_write.name());
      $display("gen_write_strobes : 'b%b", gen_write_strobes );
      $display("operation_mode   : %s", operation_mode.name() );
      $display("delay_mode       : %s", delay_mode.name() );
      $display("write_data_mode  : %s", write_data_mode.name() );
      foreach( data_beat_done[i0_1] )
        $display("data_beat_done[%0d] : 'b%b", i0_1, data_beat_done[i0_1] );
      $display("transaction_done : 'b%b", transaction_done );
      if ( print_delays == 1'b1 )
      begin
        $display("address_valid_delay : %0d", address_valid_delay);
        foreach( data_valid_delay[i0_1] )
          $display("data_valid_delay[%0d] : %0d", i0_1, data_valid_delay[i0_1]);
        $display("write_response_valid_delay : %0d", write_response_valid_delay);
        $display("address_ready_delay : %0d", address_ready_delay);
        foreach( data_ready_delay[i0_1] )
          $display("data_ready_delay[%0d] : %0d", i0_1, data_ready_delay[i0_1]);
        $display("write_response_ready_delay : %0d", write_response_ready_delay);
      end
    endfunction
endclass

`endif // MODEL_TECH
endpackage

import mgc_axi_pkg::*;
`ifdef MODEL_TECH
// *****************************************************************************
//
// Copyright 2007-2016 Mentor Graphics Corporation
// All Rights Reserved.
//
// THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE PROPERTY OF
// MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS.
//
// *****************************************************************************
// SystemVerilog           Version: 20160107
// *****************************************************************************

import QUESTA_MVC::questa_mvc_reporter;
import QUESTA_MVC::questa_mvc_item_comms_semantic;
import QUESTA_MVC::questa_mvc_edge;
import QUESTA_MVC::QUESTA_MVC_POSEDGE;
import QUESTA_MVC::QUESTA_MVC_NEGEDGE;
import QUESTA_MVC::QUESTA_MVC_ANYEDGE;
import QUESTA_MVC::QUESTA_MVC_0_TO_1_EDGE;
import QUESTA_MVC::QUESTA_MVC_1_TO_0_EDGE;


(* cy_so="libaxi_IN_SystemVerilog_MTI_full" *)
(* on_lib_load="axi_IN_SystemVerilog_load" *)

interface mgc_common_axi #(int AXI_ADDRESS_WIDTH = 64, int AXI_RDATA_WIDTH = 1024, int AXI_WDATA_WIDTH = 1024, int AXI_ID_WIDTH = 18)
    (input wire iACLK, input wire iARESETn);

    //-------------------------------------------------------------------------
    //
    // Group: AXI Signals
    //
    //-------------------------------------------------------------------------



    //-------------------------------------------------------------------------
    // Private wires
    //-------------------------------------------------------------------------
    wire ACLK;
    wire ARESETn;
    wire AWVALID;
    wire [((AXI_ADDRESS_WIDTH) - 1):0]  AWADDR;
    wire [3:0] AWLEN;
    wire [2:0] AWSIZE;
    wire [1:0] AWBURST;
    wire [1:0] AWLOCK;
    wire [3:0] AWCACHE;
    wire [2:0] AWPROT;
    wire [((AXI_ID_WIDTH) - 1):0]  AWID;
    wire AWREADY;
    wire [7:0] AWUSER;
    wire ARVALID;
    wire [((AXI_ADDRESS_WIDTH) - 1):0]  ARADDR;
    wire [3:0] ARLEN;
    wire [2:0] ARSIZE;
    wire [1:0] ARBURST;
    wire [1:0] ARLOCK;
    wire [3:0] ARCACHE;
    wire [2:0] ARPROT;
    wire [((AXI_ID_WIDTH) - 1):0]  ARID;
    wire ARREADY;
    wire [7:0] ARUSER;
    wire RVALID;
    wire RLAST;
    wire [((AXI_RDATA_WIDTH) - 1):0]  RDATA;
    wire [1:0] RRESP;
    wire [((AXI_ID_WIDTH) - 1):0]  RID;
    wire RREADY;
    wire [7:0] RUSER;
    wire WVALID;
    wire WLAST;
    wire [((AXI_WDATA_WIDTH) - 1):0]  WDATA;
    wire [(((AXI_WDATA_WIDTH / 8)) - 1):0]  WSTRB;
    wire [((AXI_ID_WIDTH) - 1):0]  WID;
    wire WREADY;
    wire [7:0] WUSER;
    wire BVALID;
    wire [1:0] BRESP;
    wire [((AXI_ID_WIDTH) - 1):0]  BID;
    wire BREADY;
    wire [7:0] BUSER;



    // Propagate global signals onto interface wires
    assign ACLK = iACLK;
    assign ARESETn = iARESETn;

    // Variable: config_write_ctrl_to_data_mintime
    //
    // 
    // Sets the delay from start of address phase to start of data phase in a write 
    // transaction (in terms of ACLK).
    // 
    // Default: 1 
    // 
    // This configuration variable has been deprecated and is maintained 
    // for backward compatibility. However, you can use ~write_address_to_data_delay~ 
    // configuration variable to control the delay between a write address phase 
    // and a write data phase.
    // 
    //
    int unsigned config_write_ctrl_to_data_mintime;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Enables
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_enable_all_assertions
    //
    // 
    // Enables all protocol assertions. 
    // 
    // Default: 1
    // 
    //
    // mentor configurator specification name "Enable all protocol assertions"
    bit config_enable_all_assertions;

    // Variable: config_enable_assertion
    //
    // 
    // Enables individual protocol assertion.
    // This variable controls whether specific assertion within QVIP (of type <axi_assertion_e>) is enabled or disabled.
    // Individual assertion can be disabled as follows:-
    // //-----------------------------------------------------------------------
    // // < BFM interface>.set_config_enable_assertion_index1(<name of assertion>,1'b0);
    // //-----------------------------------------------------------------------
    // 
    // For example, the assertion AXI_READ_DATA_UNKN is disabled as follows:
    // <bfm>.set_config_enable_assertion_index1(AXI_READ_DATA_UNKN, 1'b0); 
    // 
    // Here bfm is the AXI interface instance name for which the assertion to be disabled. 
    // 
    // Default: All assertions are enabled
    //   
    // 
    //
    // mentor configurator specification name "Enable individual protocol assertion"
    bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Slave behavior control
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_support_exclusive_access
    //
    // 
    // Enables exclusive transactions support for slave.
    // If disabled, every exclusive read/write returns an OKAY response,
    // and exclusive write updates memory. 
    // 
    // Default: 1  
    // 
    //
    // mentor configurator specification name "Enable exclusive transaction support"
    bit config_support_exclusive_access;

    // Variable: config_read_data_reordering_depth
    //
    // 
    // Sets the maximum number of different read transaction addresses for which read 
    // data(response) can be sent in any order from slave. 
    // 
    // Default: 2 ** AXI_ID_WIDTH
    // 
    //
    // mentor configurator specification name "Read data reordering depth"
    int unsigned config_read_data_reordering_depth;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Timeout control
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_max_transaction_time_factor
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) for any complete read or write transaction, which
    // includes time period for all individual phases of transaction. 
    // 
    // Default: 100000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout for complete read/write transaction"
    int unsigned config_max_transaction_time_factor;

    // Variable: config_timeout_max_data_transfer
    //
    //  
    // Sets maximum number of write data beats in a write data burst. 
    // 
    // Default: 1024  
    // 
    //
    // mentor configurator specification name "Maximum number of data beats in a write data burst"
    int config_timeout_max_data_transfer;

    // Variable: config_burst_timeout_factor
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) between individual phases of a transaction. 
    // 
    // Default: 10000 clock cycles 
    // 
    //
    // mentor configurator specification name "Burst timeout between individual phases of a transaction"
    int unsigned config_burst_timeout_factor;

    // Variable: config_max_latency_AWVALID_assertion_to_AWREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of AWVALID to assertion of AWREADY.
    // An error message AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID is generated if AWREADY is not asserted
    // after assertion of AWVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from AWVALID to AWREADY assertion"
    int unsigned config_max_latency_AWVALID_assertion_to_AWREADY;

    // Variable: config_max_latency_ARVALID_assertion_to_ARREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of ARVALID to assertion of ARREADY.
    // An error message AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID is generated if ARREADY is not asserted
    // after assertion of ARVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from ARVALID to ARREADY assertion"
    int unsigned config_max_latency_ARVALID_assertion_to_ARREADY;

    // Variable: config_max_latency_RVALID_assertion_to_RREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of RVALID to assertion of RREADY.
    // An error message AXI_RREADY_NOT_ASSERTED_AFTER_RVALID is generated if RREADY is not asserted
    // after assertion of RVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from RVALID to RREADY assertion"
    int unsigned config_max_latency_RVALID_assertion_to_RREADY;

    // Variable: config_max_latency_BVALID_assertion_to_BREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of BVALID to assertion of BREADY.
    // An error message AXI_BREADY_NOT_ASSERTED_AFTER_BVALID is generated if BREADY is not asserted
    // after assertion of BVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from BVALID to BREADY assertion"
    int unsigned config_max_latency_BVALID_assertion_to_BREADY;

    // Variable: config_max_latency_WVALID_assertion_to_WREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of WVALID to assertion of WREADY.
    // An error message AXI_WREADY_NOT_ASSERTED_AFTER_WVALID is generated if WREADY is not asserted
    // after assertion of WVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from WVALID to WREADY assertion"
    int unsigned config_max_latency_WVALID_assertion_to_WREADY;

    // Variable: config_setup_time
    //
    // 
    // Sets number of simulation time units from the setup time to the active 
    // clock edge of ACLK. The setup time will always be less than the time period
    // of the clock. 
    // 
    // Default: 0
    // 
    //
    // Note - This configuration variable is used in an expression involving time precision.
    //        To ensure its value is correct, use questa_mvc_sv_convert_to_precision API of QUESTA_MVC package.
    //
    int config_setup_time;

    // Variable: config_hold_time
    //
    // 
    // Sets number of simulation time units from the hold time to the active 
    // clock edge of ACLK. 
    // 
    // Default: 0
    // 
    //
    // Note - This configuration variable is used in an expression involving time precision.
    //        To ensure its value is correct, use questa_mvc_sv_convert_to_precision API of QUESTA_MVC package.
    //
    int config_hold_time;

    // Variable: config_max_outstanding_wr
    //
    // Configures maximum possible outstanding Write transactions
    //
    int config_max_outstanding_wr;

    // Variable: config_max_outstanding_rd
    //
    // Configures maximum possible outstanding Read transactions
    //
    int config_max_outstanding_rd;

    // Variable: config_max_outstanding_rw
    //
    // Configures maximum possible outstanding Combined (Read and Write) transactions
    //
    int config_max_outstanding_rw;

    // Variable: config_is_issuing
    //
    // Enables Master component to use "config_max_outstanding_wr/config_max_outstanding_rd/config_max_outstanding_rw" variables for transaction issuing capability when set to true
    //
    bit config_is_issuing;


    //-------------------------------------------------------------------------
    // Deprecated variables - writing to these variables will cause a warning to be issued.
    //-------------------------------------------------------------------------
    bit config_master_write_delay;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr;
    axi_error_e config_master_error_position;
    //------------------------------------------------------------------------------
    // Group:- Interface ends
    //------------------------------------------------------------------------------
    //
    longint axi_master_end;


    // Function:- get_axi_master_end
    //
    // Returns a handle to the <master> end of this instance of the <axi> interface.

    function longint get_axi_master_end();
        return axi_master_end;
    endfunction

    longint axi_slave_end;


    // Function:- get_axi_slave_end
    //
    // Returns a handle to the <slave> end of this instance of the <axi> interface.

    function longint get_axi_slave_end();
        return axi_slave_end;
    endfunction

    longint axi_clock_source_end;


    // Function:- get_axi_clock_source_end
    //
    // Returns a handle to the <clock_source> end of this instance of the <axi> interface.

    function longint get_axi_clock_source_end();
        return axi_clock_source_end;
    endfunction

    longint axi_reset_source_end;


    // Function:- get_axi_reset_source_end
    //
    // Returns a handle to the <reset_source> end of this instance of the <axi> interface.

    function longint get_axi_reset_source_end();
        return axi_reset_source_end;
    endfunction

    longint axi__monitor_end;


    // Function:- get_axi__monitor_end
    //
    // Returns a handle to the <_monitor> end of this instance of the <axi> interface.

    function longint get_axi__monitor_end();
        return axi__monitor_end;
    endfunction


    // Group:- Abstraction Levels
    // 
    // These functions are used set or get the abstraction levels of an interface end.
    // See <Abstraction Levels of Interface Ends> for more details on the meaning of
    // TLM or WLM connected and the valid combinations.


    //-------------------------------------------------------------------------
    // Function:- axi_set_master_abstraction_level
    //
    //     Function to set whether the <master> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_master_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_master_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_master_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <master> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_master_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_master_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_slave_abstraction_level
    //
    //     Function to set whether the <slave> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_slave_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_slave_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_slave_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <slave> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_slave_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_slave_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_clock_source_abstraction_level
    //
    //     Function to set whether the <clock_source> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_clock_source_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_clock_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_clock_source_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <clock_source> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_clock_source_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_clock_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_reset_source_abstraction_level
    //
    //     Function to set whether the <reset_source> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_reset_source_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_reset_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_reset_source_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <reset_source> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_reset_source_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_reset_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    import "DPI-C" context function longint axi_initialise_SystemVerilog
    (
        int    usage_code,
        string iface_version,
        output longint master_end,
        output longint slave_end,
        output longint clock_source_end,
        output longint reset_source_end,
        output longint _monitor_end,
        input int AXI_ADDRESS_WIDTH,
        input int AXI_RDATA_WIDTH,
        input int AXI_WDATA_WIDTH,
        input int AXI_ID_WIDTH
    );

    `ifndef MVC_axi_VERSION
    `define MVC_axi_VERSION ""
    `endif
    // Handle to the linkage
    (* elab_init *) longint _interface_ref =
                                axi_initialise_SystemVerilog
                                (
                                    18102076,
                                    `MVC_axi_VERSION,
                                    axi_master_end,
                                    axi_slave_end,
                                    axi_clock_source_end,
                                    axi_reset_source_end,
                                    axi__monitor_end,
                                    AXI_ADDRESS_WIDTH,
                                    AXI_RDATA_WIDTH,
                                    AXI_WDATA_WIDTH,
                                    AXI_ID_WIDTH
                                ); // DPI call to create transactor (called at
                                     // elaboration time as initialiser)

    generate
    begin : questa_mvc_reporting
        bit report_available;

        // Function for getting a message from QUESTA_MVC. Returns 1 if a message was returned, 0 otherwise.
        import "DPI-C" questa_mvc_sv_get_report =  function bit get_report( input longint iface_ref,input longint recipient,
                                     output string category,     output string objectName,
                                     output string instanceName, output string error_no,
                                     output string typ,          output string mess );
        questa_mvc_reporter endPoint[longint];
        initial report_available = 0;

        always @report_available
        begin
            longint recipient;
            string category;
            string objectName;
            string instanceName;
            string severity;
            string mess;
            string error_no;

            if ( endPoint.first( recipient ) )
              begin
                do
                  begin
                      while ( get_report( _interface_ref, recipient, category, objectName, instanceName, error_no, severity, mess ) )
                        begin
                          endPoint[recipient].report_message( category, "axi", 0, objectName, instanceName, error_no, severity, mess );
                        end
                  end
                while (endPoint.next(recipient));
              end
            report_available = 0;
        end

        import "DPI-C" context questa_mvc_register_end_point = function void questa_mvc_register_end_point( input longint iface_ref, input longint as_end, input string name );

        // A function for registering a reporter to capture any reports coming from as_end
        function automatic void register_end_point( input longint as_end, input questa_mvc_reporter rep = null );
            if ( rep != null )
              begin
                if ( ( rep.name == "" ) || ( rep.name == "NULL" ) )
                  begin
                    $display("Error: %m: Reporter passed to register_end_point has a reserved name. Neither an empty string nor the string 'NULL' can be used.");
                  end
                else
                  begin
                    questa_mvc_register_end_point( _interface_ref, as_end, rep.name );
                    endPoint[as_end] = rep;
                  end
              end
            else
              begin
                questa_mvc_register_end_point( _interface_ref, as_end, "NULL" );
                endPoint.delete( as_end );
              end
        endfunction

    end : questa_mvc_reporting
    endgenerate

    //-------------------------------------------------------------------------
    //
    // Group:- Registering Reports
    //
    //
    // The following methods are used to register a custom reporting object as
    // described in the MVC base library section, <Customizing Error-Reporting>.
    // 
    //-------------------------------------------------------------------------

    function void register_interface_reporter( input questa_mvc_reporter _rep = null );
        questa_mvc_reporting.register_end_point( _interface_ref, _rep );
    endfunction


    // Support the old API for registering an interface, for backwards compatability.
    // Note that this function is deprecated and may be removed in the future.
    function void interface_register_reporter( input questa_mvc_reporter _rep = null );
        questa_mvc_reporting.register_end_point( _interface_ref, _rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_master_reporter
    //
    // Function used to register a reporter for the <master> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the master end.
    //
    function void register_master_reporter
    (
        input questa_mvc_reporter rep = null
    );
        questa_mvc_reporting.register_end_point( axi_master_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_slave_reporter
    //
    // Function used to register a reporter for the <slave> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the slave end.
    //
    function void register_slave_reporter
    (
        input questa_mvc_reporter rep = null
    );
        questa_mvc_reporting.register_end_point( axi_slave_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_clock_source_reporter
    //
    // Function used to register a reporter for the <clock_source> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the clock_source end.
    //
    function void register_clock_source_reporter
    (
        input questa_mvc_reporter rep = null
    );
        questa_mvc_reporting.register_end_point( axi_clock_source_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_reset_source_reporter
    //
    // Function used to register a reporter for the <reset_source> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the reset_source end.
    //
    function void register_reset_source_reporter
    (
        input questa_mvc_reporter rep = null
    );
        questa_mvc_reporting.register_end_point( axi_reset_source_end, rep );
    endfunction


    //-------------------------------------------------------------------------
    //
    // Group: BFM Utility/Convenience Methods
    //
    // This is the group of utility functions provided by the QVIP BFM to
    // communicate from the SV world to the QVIP BFM.
    // This set of APIs can be used to either get status/statistics
    // information from the BFM or to set values in a particular database 
    // in the BFM. Please refer to individual functions for more information.
    //
    //-------------------------------------------------------------------------

    //-------------------------------------------------------------------------
    // Function: fn_rd_txn_valid_lanes
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get valid strobes/lanes value for each of the read data beat
    //     at end of read transaction.
    // 
    //     Please note that this function should be called after completion of a read
    //     transaction.
    // 
    //     Output of the function:
    //     valid_lanes - Valid strobes value for each read data beat
    //    
    function automatic void fn_rd_txn_valid_lanes
    (
        ref bit [((AXI_RDATA_WIDTH / 8) - 1):0] valid_lanes []
    );
         fn_rd_txn_valid_lanes_C(valid_lanes);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_get_wdata_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get information corresponding to a write data beat.
    // 
    //     Input:
    //     id         - ID of the write data beat
    //     wdata_last - assigned to ~last~ attribute of the write data beat
    // 
    //     Output:
    //     waddr_rcvd   - Indicates if corresponding write address phase is received
    //     burst_length - Burst length attribute of the corresponding address phase
    //     beat_num     - Write data beat number of the corresponding write data burst
    //     beat_addr    - Corresponding beat address
    // 
    //     Please note that this function should be called at the completion of write
    //     data beat.
    //    
    function automatic void fn_get_wdata_phase_info
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit wdata_last,
        inout bit waddr_rcvd,
        output bit [3:0] burst_length,
        output int beat_num,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  beat_addr
    );
         fn_get_wdata_phase_info_C(id,wdata_last,waddr_rcvd,burst_length,beat_num,beat_addr);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_get_wresp_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get address attribute of write address phase corresponding
    //     to write response phase that just completed.
    // 
    //     Please note that this function should be called after completion of a write
    //     response phase.
    // 
    //     Output of the function:
    //     wresp_corr_addr - ~addr~ attribute of the address phase corresponding to
    //                       this write response phase
    //    
    function automatic void fn_get_wresp_phase_info
    (
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  wresp_corr_addr
    );
         fn_get_wresp_phase_info_C(wresp_corr_addr);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_get_rdata_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get information corresponding to a read data beat.
    // 
    //     Input:
    //     id         - ID of the read data beat
    // 
    //     Output:
    //     burst_length - Burst length attribute of the corresponding read address phase
    //     beat_num     - Read data beat number of the corresponding read data burst
    //     beat_strobes - Valid lanes in the read data beat
    //     beat_addr    - Corresponding beat address
    // 
    //     Please note that this function should be called at the completion of read
    //     data beat.
    //    
    function automatic void fn_get_rdata_phase_info
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit rdata_last,
        output bit [3:0] burst_length,
        output int beat_num,
        output bit [((AXI_RDATA_WIDTH / 8) - 1):0]  beat_strobes,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  beat_addr,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  txn_addr
    );
         fn_get_rdata_phase_info_C(id,rdata_last,burst_length,beat_num,beat_strobes,beat_addr,txn_addr);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_get_max_os_per_id
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function gets the maximum number of outstanding write phases of a particular ID
    // from among all AWID, WID values.
    //  
    // Inputs:
    // max_waddr_os - The maximum number of address phases outstanding from among all AWID
    // max_wdata_os - The maximum number of data bursts outstanding from among all WID
    // 
    // For example, 5 write address phases are outstanding with ID 3, and 
    // 7 write address phases are outstanding with ID 2. No other address phase is there
    // and 0 write data phases are received.
    // 
    // The return values would be such that:
    // max_waddr_os = 7
    // max_wdata_os = 0
    // 
    function automatic void fn_get_max_os_per_id
    (
        output int max_waddr_os,
        output int max_wdata_os
    );
         fn_get_max_os_per_id_C(max_waddr_os,max_wdata_os);
    endfunction

    //-------------------------------------------------------------------------
    // Function: get_rw_txns_in_prog
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function gets the number of various outstanding transactions at a time.
    // 
    // Inputs:
    // id  - The AWID/ARID/WID of the transaction whose details are required.
    // txn_counts - The statistics of the number of outstanding transactions
    function automatic void get_rw_txns_in_prog
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_rw_txn_counts_s txn_counts
    );
         get_rw_txns_in_prog_C(id,txn_counts);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_add_addr_map_entry
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets address map fields inside internal BFM. 
    // 
    // Inputs:
    // region - Region name 
    // addr - Start address of region
    // size - Size of address region
    function automatic void fn_add_addr_map_entry
    (
        input string region,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input longint unsigned size
    );
         fn_add_addr_map_entry_C(region,addr,size);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_add_wr_delay
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets delay values for write address-data pair and 
    // between write data beats, initiated by master end. 
    // 
    // Inputs:
    // region - Region value for which write delays are to be inserted
    // id - Write transaction's id (AWID) for which delays are to be inserted
    // addr2data - Delays to be inserted between write address and data phase.
    // data2data - Delays to be inserted between data beats
    function automatic void fn_add_wr_delay
    (
        input string region,
        input bit [17:0] id,
        input int unsigned addr2data,
        ref int unsigned data2data[]
    );
         fn_add_wr_delay_C(region,id,addr2data,data2data);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_delete_wr_delay
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function deletes delay values for a region-id pair
    // 
    // Inputs:
    // region - Region value for which write delays are to be inserted
    // id - Write transaction's id (AWID) for which delays are to be inserted
    // addr2data - Delays to be inserted between write address and data phase.
    // data2data - Delays to be inserted between data beats
    function automatic void fn_delete_wr_delay
    (
        input string region,
        input bit [17:0] id
    );
         fn_delete_wr_delay_C(region,id);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_set_wr_def_delays
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets default delay values for write address-data pair and data beats 
    // initiated by master end between input max. and min. values. In case non-randomized 
    // default value is desired, user can set max. and min. to same value.
    // 
    // Inputs:
    // min_addr2data - Minimum value of default delays to be inserted between write address and data phase.
    // min_data2data - Minimum value of default delays to be inserted between data beats
    // max_addr2data - Maximum value of default delays to be inserted between write address and data phase.
    // max_data2data - Maximum value of default delays to be inserted between data beats
    function automatic void fn_set_wr_def_delays
    (
        input int unsigned min_addr2data,
        ref int unsigned min_data2data[],
        input int unsigned max_addr2data,
        ref int unsigned max_data2data[]
    );
         fn_set_wr_def_delays_C(min_addr2data,min_data2data,max_addr2data,max_data2data);
    endfunction

    // Declare user visible wires variables, for non-continuous assignments.
    logic m_ACLK = 'z;
    logic m_ARESETn = 'z;
    logic m_AWVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  m_AWADDR = 'z;
    logic [3:0] m_AWLEN = 'z;
    logic [2:0] m_AWSIZE = 'z;
    logic [1:0] m_AWBURST = 'z;
    logic [1:0] m_AWLOCK = 'z;
    logic [3:0] m_AWCACHE = 'z;
    logic [2:0] m_AWPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_AWID = 'z;
    logic m_AWREADY = 'z;
    logic [7:0] m_AWUSER = 'z;
    logic m_ARVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  m_ARADDR = 'z;
    logic [3:0] m_ARLEN = 'z;
    logic [2:0] m_ARSIZE = 'z;
    logic [1:0] m_ARBURST = 'z;
    logic [1:0] m_ARLOCK = 'z;
    logic [3:0] m_ARCACHE = 'z;
    logic [2:0] m_ARPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_ARID = 'z;
    logic m_ARREADY = 'z;
    logic [7:0] m_ARUSER = 'z;
    logic m_RVALID = 'z;
    logic m_RLAST = 'z;
    logic [((AXI_RDATA_WIDTH) - 1):0]  m_RDATA = 'z;
    logic [1:0] m_RRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_RID = 'z;
    logic m_RREADY = 'z;
    logic [7:0] m_RUSER = 'z;
    logic m_WVALID = 'z;
    logic m_WLAST = 'z;
    logic [((AXI_WDATA_WIDTH) - 1):0]  m_WDATA = 'z;
    logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  m_WSTRB = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_WID = 'z;
    logic m_WREADY = 'z;
    logic [7:0] m_WUSER = 'z;
    logic m_BVALID = 'z;
    logic [1:0] m_BRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_BID = 'z;
    logic m_BREADY = 'z;
    logic [7:0] m_BUSER = 'z;

    // Forces a sweep through the wire change checkers at time 0 to get around
    // process kick-off order unknowns
    bit _check_t0_values;
    always_comb _check_t0_values = 1;

    // handle control
    longint last_handle = 0;

    longint last_start_time = 0;

    longint last_end_time = 0;

    export "DPI-C" axi_set_last_handle_and_times = function set_last_handle_and_times;

    function void set_last_handle_and_times(longint _handle, longint _start, longint _end);
        last_handle = _handle;
        last_start_time = _start;
        last_end_time = _end;
    endfunction


    function longint get_last_handle();
        return last_handle;
    endfunction


    function longint get_last_start_time();
        return last_start_time;
    endfunction


    function longint get_last_end_time();
        return last_end_time;
    endfunction


    //-------------------------------------------------------------------------
    // Tasks to wait for a number of specified edges on a wire
    //-------------------------------------------------------------------------


    //------------------------------------------------------------------------------
    // Function:- wait_for_ACLK
    //     Wait for the specified change on wire <axi::ACLK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ACLK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ACLK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ACLK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ACLK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ACLK === 0 );
                    @( ACLK );
                end
                while ( ACLK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ACLK === 1 );
                    @( ACLK );
                end
                while ( ACLK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARESETn
    //     Wait for the specified change on wire <axi::ARESETn>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARESETn( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARESETn);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARESETn);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARESETn);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARESETn === 0 );
                    @( ARESETn );
                end
                while ( ARESETn !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARESETn === 1 );
                    @( ARESETn );
                end
                while ( ARESETn !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWVALID
    //     Wait for the specified change on wire <axi::AWVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWVALID === 0 );
                    @( AWVALID );
                end
                while ( AWVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWVALID === 1 );
                    @( AWVALID );
                end
                while ( AWVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWADDR
    //     Wait for the specified change on wire <axi::AWADDR>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWADDR( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWADDR);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWADDR);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWADDR);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWADDR === 0 );
                    @( AWADDR );
                end
                while ( AWADDR !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWADDR === 1 );
                    @( AWADDR );
                end
                while ( AWADDR !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWADDR_index1
    //     Wait for the specified change on wire <axi::AWADDR>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWADDR_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWADDR[_this_dot_1] === 0 );
                    @( AWADDR[_this_dot_1] );
                end
                while ( AWADDR[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWADDR[_this_dot_1] === 1 );
                    @( AWADDR[_this_dot_1] );
                end
                while ( AWADDR[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLEN
    //     Wait for the specified change on wire <axi::AWLEN>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLEN( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLEN);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLEN);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLEN);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLEN === 0 );
                    @( AWLEN );
                end
                while ( AWLEN !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLEN === 1 );
                    @( AWLEN );
                end
                while ( AWLEN !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLEN_index1
    //     Wait for the specified change on wire <axi::AWLEN>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLEN_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLEN[_this_dot_1] === 0 );
                    @( AWLEN[_this_dot_1] );
                end
                while ( AWLEN[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLEN[_this_dot_1] === 1 );
                    @( AWLEN[_this_dot_1] );
                end
                while ( AWLEN[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWSIZE
    //     Wait for the specified change on wire <axi::AWSIZE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWSIZE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWSIZE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWSIZE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWSIZE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWSIZE === 0 );
                    @( AWSIZE );
                end
                while ( AWSIZE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWSIZE === 1 );
                    @( AWSIZE );
                end
                while ( AWSIZE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWSIZE_index1
    //     Wait for the specified change on wire <axi::AWSIZE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWSIZE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWSIZE[_this_dot_1] === 0 );
                    @( AWSIZE[_this_dot_1] );
                end
                while ( AWSIZE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWSIZE[_this_dot_1] === 1 );
                    @( AWSIZE[_this_dot_1] );
                end
                while ( AWSIZE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWBURST
    //     Wait for the specified change on wire <axi::AWBURST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWBURST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWBURST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWBURST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWBURST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWBURST === 0 );
                    @( AWBURST );
                end
                while ( AWBURST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWBURST === 1 );
                    @( AWBURST );
                end
                while ( AWBURST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWBURST_index1
    //     Wait for the specified change on wire <axi::AWBURST>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWBURST_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWBURST[_this_dot_1] === 0 );
                    @( AWBURST[_this_dot_1] );
                end
                while ( AWBURST[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWBURST[_this_dot_1] === 1 );
                    @( AWBURST[_this_dot_1] );
                end
                while ( AWBURST[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLOCK
    //     Wait for the specified change on wire <axi::AWLOCK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLOCK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLOCK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLOCK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLOCK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLOCK === 0 );
                    @( AWLOCK );
                end
                while ( AWLOCK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLOCK === 1 );
                    @( AWLOCK );
                end
                while ( AWLOCK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLOCK_index1
    //     Wait for the specified change on wire <axi::AWLOCK>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLOCK_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLOCK[_this_dot_1] === 0 );
                    @( AWLOCK[_this_dot_1] );
                end
                while ( AWLOCK[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLOCK[_this_dot_1] === 1 );
                    @( AWLOCK[_this_dot_1] );
                end
                while ( AWLOCK[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWCACHE
    //     Wait for the specified change on wire <axi::AWCACHE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWCACHE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWCACHE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWCACHE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWCACHE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWCACHE === 0 );
                    @( AWCACHE );
                end
                while ( AWCACHE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWCACHE === 1 );
                    @( AWCACHE );
                end
                while ( AWCACHE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWCACHE_index1
    //     Wait for the specified change on wire <axi::AWCACHE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWCACHE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWCACHE[_this_dot_1] === 0 );
                    @( AWCACHE[_this_dot_1] );
                end
                while ( AWCACHE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWCACHE[_this_dot_1] === 1 );
                    @( AWCACHE[_this_dot_1] );
                end
                while ( AWCACHE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWPROT
    //     Wait for the specified change on wire <axi::AWPROT>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWPROT( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWPROT);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWPROT);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWPROT);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWPROT === 0 );
                    @( AWPROT );
                end
                while ( AWPROT !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWPROT === 1 );
                    @( AWPROT );
                end
                while ( AWPROT !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWPROT_index1
    //     Wait for the specified change on wire <axi::AWPROT>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWPROT_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWPROT[_this_dot_1] === 0 );
                    @( AWPROT[_this_dot_1] );
                end
                while ( AWPROT[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWPROT[_this_dot_1] === 1 );
                    @( AWPROT[_this_dot_1] );
                end
                while ( AWPROT[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWID
    //     Wait for the specified change on wire <axi::AWID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWID === 0 );
                    @( AWID );
                end
                while ( AWID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWID === 1 );
                    @( AWID );
                end
                while ( AWID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWID_index1
    //     Wait for the specified change on wire <axi::AWID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWID[_this_dot_1] === 0 );
                    @( AWID[_this_dot_1] );
                end
                while ( AWID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWID[_this_dot_1] === 1 );
                    @( AWID[_this_dot_1] );
                end
                while ( AWID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWREADY
    //     Wait for the specified change on wire <axi::AWREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWREADY === 0 );
                    @( AWREADY );
                end
                while ( AWREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWREADY === 1 );
                    @( AWREADY );
                end
                while ( AWREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWUSER
    //     Wait for the specified change on wire <axi::AWUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWUSER === 0 );
                    @( AWUSER );
                end
                while ( AWUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWUSER === 1 );
                    @( AWUSER );
                end
                while ( AWUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWUSER_index1
    //     Wait for the specified change on wire <axi::AWUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWUSER[_this_dot_1] === 0 );
                    @( AWUSER[_this_dot_1] );
                end
                while ( AWUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWUSER[_this_dot_1] === 1 );
                    @( AWUSER[_this_dot_1] );
                end
                while ( AWUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARVALID
    //     Wait for the specified change on wire <axi::ARVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARVALID === 0 );
                    @( ARVALID );
                end
                while ( ARVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARVALID === 1 );
                    @( ARVALID );
                end
                while ( ARVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARADDR
    //     Wait for the specified change on wire <axi::ARADDR>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARADDR( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARADDR);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARADDR);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARADDR);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARADDR === 0 );
                    @( ARADDR );
                end
                while ( ARADDR !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARADDR === 1 );
                    @( ARADDR );
                end
                while ( ARADDR !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARADDR_index1
    //     Wait for the specified change on wire <axi::ARADDR>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARADDR_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARADDR[_this_dot_1] === 0 );
                    @( ARADDR[_this_dot_1] );
                end
                while ( ARADDR[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARADDR[_this_dot_1] === 1 );
                    @( ARADDR[_this_dot_1] );
                end
                while ( ARADDR[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLEN
    //     Wait for the specified change on wire <axi::ARLEN>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLEN( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLEN);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLEN);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLEN);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLEN === 0 );
                    @( ARLEN );
                end
                while ( ARLEN !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLEN === 1 );
                    @( ARLEN );
                end
                while ( ARLEN !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLEN_index1
    //     Wait for the specified change on wire <axi::ARLEN>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLEN_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLEN[_this_dot_1] === 0 );
                    @( ARLEN[_this_dot_1] );
                end
                while ( ARLEN[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLEN[_this_dot_1] === 1 );
                    @( ARLEN[_this_dot_1] );
                end
                while ( ARLEN[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARSIZE
    //     Wait for the specified change on wire <axi::ARSIZE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARSIZE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARSIZE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARSIZE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARSIZE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARSIZE === 0 );
                    @( ARSIZE );
                end
                while ( ARSIZE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARSIZE === 1 );
                    @( ARSIZE );
                end
                while ( ARSIZE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARSIZE_index1
    //     Wait for the specified change on wire <axi::ARSIZE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARSIZE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARSIZE[_this_dot_1] === 0 );
                    @( ARSIZE[_this_dot_1] );
                end
                while ( ARSIZE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARSIZE[_this_dot_1] === 1 );
                    @( ARSIZE[_this_dot_1] );
                end
                while ( ARSIZE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARBURST
    //     Wait for the specified change on wire <axi::ARBURST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARBURST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARBURST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARBURST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARBURST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARBURST === 0 );
                    @( ARBURST );
                end
                while ( ARBURST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARBURST === 1 );
                    @( ARBURST );
                end
                while ( ARBURST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARBURST_index1
    //     Wait for the specified change on wire <axi::ARBURST>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARBURST_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARBURST[_this_dot_1] === 0 );
                    @( ARBURST[_this_dot_1] );
                end
                while ( ARBURST[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARBURST[_this_dot_1] === 1 );
                    @( ARBURST[_this_dot_1] );
                end
                while ( ARBURST[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLOCK
    //     Wait for the specified change on wire <axi::ARLOCK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLOCK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLOCK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLOCK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLOCK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLOCK === 0 );
                    @( ARLOCK );
                end
                while ( ARLOCK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLOCK === 1 );
                    @( ARLOCK );
                end
                while ( ARLOCK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLOCK_index1
    //     Wait for the specified change on wire <axi::ARLOCK>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLOCK_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLOCK[_this_dot_1] === 0 );
                    @( ARLOCK[_this_dot_1] );
                end
                while ( ARLOCK[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLOCK[_this_dot_1] === 1 );
                    @( ARLOCK[_this_dot_1] );
                end
                while ( ARLOCK[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARCACHE
    //     Wait for the specified change on wire <axi::ARCACHE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARCACHE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARCACHE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARCACHE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARCACHE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARCACHE === 0 );
                    @( ARCACHE );
                end
                while ( ARCACHE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARCACHE === 1 );
                    @( ARCACHE );
                end
                while ( ARCACHE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARCACHE_index1
    //     Wait for the specified change on wire <axi::ARCACHE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARCACHE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARCACHE[_this_dot_1] === 0 );
                    @( ARCACHE[_this_dot_1] );
                end
                while ( ARCACHE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARCACHE[_this_dot_1] === 1 );
                    @( ARCACHE[_this_dot_1] );
                end
                while ( ARCACHE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARPROT
    //     Wait for the specified change on wire <axi::ARPROT>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARPROT( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARPROT);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARPROT);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARPROT);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARPROT === 0 );
                    @( ARPROT );
                end
                while ( ARPROT !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARPROT === 1 );
                    @( ARPROT );
                end
                while ( ARPROT !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARPROT_index1
    //     Wait for the specified change on wire <axi::ARPROT>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARPROT_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARPROT[_this_dot_1] === 0 );
                    @( ARPROT[_this_dot_1] );
                end
                while ( ARPROT[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARPROT[_this_dot_1] === 1 );
                    @( ARPROT[_this_dot_1] );
                end
                while ( ARPROT[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARID
    //     Wait for the specified change on wire <axi::ARID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARID === 0 );
                    @( ARID );
                end
                while ( ARID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARID === 1 );
                    @( ARID );
                end
                while ( ARID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARID_index1
    //     Wait for the specified change on wire <axi::ARID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARID[_this_dot_1] === 0 );
                    @( ARID[_this_dot_1] );
                end
                while ( ARID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARID[_this_dot_1] === 1 );
                    @( ARID[_this_dot_1] );
                end
                while ( ARID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARREADY
    //     Wait for the specified change on wire <axi::ARREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARREADY === 0 );
                    @( ARREADY );
                end
                while ( ARREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARREADY === 1 );
                    @( ARREADY );
                end
                while ( ARREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARUSER
    //     Wait for the specified change on wire <axi::ARUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARUSER === 0 );
                    @( ARUSER );
                end
                while ( ARUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARUSER === 1 );
                    @( ARUSER );
                end
                while ( ARUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARUSER_index1
    //     Wait for the specified change on wire <axi::ARUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARUSER[_this_dot_1] === 0 );
                    @( ARUSER[_this_dot_1] );
                end
                while ( ARUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARUSER[_this_dot_1] === 1 );
                    @( ARUSER[_this_dot_1] );
                end
                while ( ARUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RVALID
    //     Wait for the specified change on wire <axi::RVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RVALID === 0 );
                    @( RVALID );
                end
                while ( RVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RVALID === 1 );
                    @( RVALID );
                end
                while ( RVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RLAST
    //     Wait for the specified change on wire <axi::RLAST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RLAST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RLAST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RLAST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RLAST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RLAST === 0 );
                    @( RLAST );
                end
                while ( RLAST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RLAST === 1 );
                    @( RLAST );
                end
                while ( RLAST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RDATA
    //     Wait for the specified change on wire <axi::RDATA>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RDATA( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RDATA);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RDATA);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RDATA);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RDATA === 0 );
                    @( RDATA );
                end
                while ( RDATA !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RDATA === 1 );
                    @( RDATA );
                end
                while ( RDATA !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RDATA_index1
    //     Wait for the specified change on wire <axi::RDATA>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RDATA_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RDATA[_this_dot_1] === 0 );
                    @( RDATA[_this_dot_1] );
                end
                while ( RDATA[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RDATA[_this_dot_1] === 1 );
                    @( RDATA[_this_dot_1] );
                end
                while ( RDATA[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RRESP
    //     Wait for the specified change on wire <axi::RRESP>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RRESP( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RRESP);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RRESP);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RRESP);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RRESP === 0 );
                    @( RRESP );
                end
                while ( RRESP !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RRESP === 1 );
                    @( RRESP );
                end
                while ( RRESP !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RRESP_index1
    //     Wait for the specified change on wire <axi::RRESP>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RRESP_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RRESP[_this_dot_1] === 0 );
                    @( RRESP[_this_dot_1] );
                end
                while ( RRESP[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RRESP[_this_dot_1] === 1 );
                    @( RRESP[_this_dot_1] );
                end
                while ( RRESP[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RID
    //     Wait for the specified change on wire <axi::RID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RID === 0 );
                    @( RID );
                end
                while ( RID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RID === 1 );
                    @( RID );
                end
                while ( RID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RID_index1
    //     Wait for the specified change on wire <axi::RID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RID[_this_dot_1] === 0 );
                    @( RID[_this_dot_1] );
                end
                while ( RID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RID[_this_dot_1] === 1 );
                    @( RID[_this_dot_1] );
                end
                while ( RID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RREADY
    //     Wait for the specified change on wire <axi::RREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RREADY === 0 );
                    @( RREADY );
                end
                while ( RREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RREADY === 1 );
                    @( RREADY );
                end
                while ( RREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RUSER
    //     Wait for the specified change on wire <axi::RUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RUSER === 0 );
                    @( RUSER );
                end
                while ( RUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RUSER === 1 );
                    @( RUSER );
                end
                while ( RUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RUSER_index1
    //     Wait for the specified change on wire <axi::RUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RUSER[_this_dot_1] === 0 );
                    @( RUSER[_this_dot_1] );
                end
                while ( RUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RUSER[_this_dot_1] === 1 );
                    @( RUSER[_this_dot_1] );
                end
                while ( RUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WVALID
    //     Wait for the specified change on wire <axi::WVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WVALID === 0 );
                    @( WVALID );
                end
                while ( WVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WVALID === 1 );
                    @( WVALID );
                end
                while ( WVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WLAST
    //     Wait for the specified change on wire <axi::WLAST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WLAST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WLAST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WLAST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WLAST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WLAST === 0 );
                    @( WLAST );
                end
                while ( WLAST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WLAST === 1 );
                    @( WLAST );
                end
                while ( WLAST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WDATA
    //     Wait for the specified change on wire <axi::WDATA>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WDATA( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WDATA);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WDATA);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WDATA);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WDATA === 0 );
                    @( WDATA );
                end
                while ( WDATA !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WDATA === 1 );
                    @( WDATA );
                end
                while ( WDATA !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WDATA_index1
    //     Wait for the specified change on wire <axi::WDATA>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WDATA_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WDATA[_this_dot_1] === 0 );
                    @( WDATA[_this_dot_1] );
                end
                while ( WDATA[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WDATA[_this_dot_1] === 1 );
                    @( WDATA[_this_dot_1] );
                end
                while ( WDATA[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WSTRB
    //     Wait for the specified change on wire <axi::WSTRB>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WSTRB( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WSTRB);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WSTRB);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WSTRB);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WSTRB === 0 );
                    @( WSTRB );
                end
                while ( WSTRB !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WSTRB === 1 );
                    @( WSTRB );
                end
                while ( WSTRB !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WSTRB_index1
    //     Wait for the specified change on wire <axi::WSTRB>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WSTRB_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WSTRB[_this_dot_1] === 0 );
                    @( WSTRB[_this_dot_1] );
                end
                while ( WSTRB[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WSTRB[_this_dot_1] === 1 );
                    @( WSTRB[_this_dot_1] );
                end
                while ( WSTRB[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WID
    //     Wait for the specified change on wire <axi::WID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WID === 0 );
                    @( WID );
                end
                while ( WID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WID === 1 );
                    @( WID );
                end
                while ( WID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WID_index1
    //     Wait for the specified change on wire <axi::WID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WID[_this_dot_1] === 0 );
                    @( WID[_this_dot_1] );
                end
                while ( WID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WID[_this_dot_1] === 1 );
                    @( WID[_this_dot_1] );
                end
                while ( WID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WREADY
    //     Wait for the specified change on wire <axi::WREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WREADY === 0 );
                    @( WREADY );
                end
                while ( WREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WREADY === 1 );
                    @( WREADY );
                end
                while ( WREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WUSER
    //     Wait for the specified change on wire <axi::WUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WUSER === 0 );
                    @( WUSER );
                end
                while ( WUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WUSER === 1 );
                    @( WUSER );
                end
                while ( WUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WUSER_index1
    //     Wait for the specified change on wire <axi::WUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WUSER[_this_dot_1] === 0 );
                    @( WUSER[_this_dot_1] );
                end
                while ( WUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WUSER[_this_dot_1] === 1 );
                    @( WUSER[_this_dot_1] );
                end
                while ( WUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BVALID
    //     Wait for the specified change on wire <axi::BVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BVALID === 0 );
                    @( BVALID );
                end
                while ( BVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BVALID === 1 );
                    @( BVALID );
                end
                while ( BVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BRESP
    //     Wait for the specified change on wire <axi::BRESP>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BRESP( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BRESP);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BRESP);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BRESP);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BRESP === 0 );
                    @( BRESP );
                end
                while ( BRESP !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BRESP === 1 );
                    @( BRESP );
                end
                while ( BRESP !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BRESP_index1
    //     Wait for the specified change on wire <axi::BRESP>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BRESP_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BRESP[_this_dot_1] === 0 );
                    @( BRESP[_this_dot_1] );
                end
                while ( BRESP[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BRESP[_this_dot_1] === 1 );
                    @( BRESP[_this_dot_1] );
                end
                while ( BRESP[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BID
    //     Wait for the specified change on wire <axi::BID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BID === 0 );
                    @( BID );
                end
                while ( BID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BID === 1 );
                    @( BID );
                end
                while ( BID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BID_index1
    //     Wait for the specified change on wire <axi::BID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BID[_this_dot_1] === 0 );
                    @( BID[_this_dot_1] );
                end
                while ( BID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BID[_this_dot_1] === 1 );
                    @( BID[_this_dot_1] );
                end
                while ( BID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BREADY
    //     Wait for the specified change on wire <axi::BREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BREADY === 0 );
                    @( BREADY );
                end
                while ( BREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BREADY === 1 );
                    @( BREADY );
                end
                while ( BREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BUSER
    //     Wait for the specified change on wire <axi::BUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BUSER === 0 );
                    @( BUSER );
                end
                while ( BUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BUSER === 1 );
                    @( BUSER );
                end
                while ( BUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BUSER_index1
    //     Wait for the specified change on wire <axi::BUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BUSER[_this_dot_1] === 0 );
                    @( BUSER[_this_dot_1] );
                end
                while ( BUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BUSER[_this_dot_1] === 1 );
                    @( BUSER[_this_dot_1] );
                end
                while ( BUSER[_this_dot_1] !== 0 );
            end
        end
    endtask

    //-------------------------------------------------------------------------
    // Tasks/functions to set/get wires
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- set_ACLK
    //-------------------------------------------------------------------------
    //     Set the value of wire <ACLK>.
    //
    // Parameters:
    //     ACLK_param - The value to set onto wire <ACLK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ACLK( logic ACLK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ACLK = ACLK_param;
        else
            m_ACLK <= ACLK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ACLK
    //-------------------------------------------------------------------------
    //     Get the value of wire <ACLK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ACLK>.
    //
    function automatic logic get_ACLK(  );
        return ACLK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARESETn
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARESETn>.
    //
    // Parameters:
    //     ARESETn_param - The value to set onto wire <ARESETn>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARESETn( logic ARESETn_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARESETn = ARESETn_param;
        else
            m_ARESETn <= ARESETn_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARESETn
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARESETn>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARESETn>.
    //
    function automatic logic get_ARESETn(  );
        return ARESETn;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWVALID>.
    //
    // Parameters:
    //     AWVALID_param - The value to set onto wire <AWVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWVALID( logic AWVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWVALID = AWVALID_param;
        else
            m_AWVALID <= AWVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWVALID>.
    //
    function automatic logic get_AWVALID(  );
        return AWVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWADDR
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWADDR>.
    //
    // Parameters:
    //     AWADDR_param - The value to set onto wire <AWADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWADDR( logic [((AXI_ADDRESS_WIDTH) - 1):0]  AWADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWADDR = AWADDR_param;
        else
            m_AWADDR <= AWADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWADDR_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWADDR_param - The value to set onto wire <AWADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWADDR_index1( int _this_dot_1, logic  AWADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWADDR[_this_dot_1] = AWADDR_param;
        else
            m_AWADDR[_this_dot_1] <= AWADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWADDR
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWADDR>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWADDR>.
    //
    function automatic logic [((AXI_ADDRESS_WIDTH) - 1):0]   get_AWADDR(  );
        return AWADDR;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWADDR_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWADDR>.
    //
    function automatic logic   get_AWADDR_index1( int _this_dot_1 );
        return AWADDR[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWLEN
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWLEN>.
    //
    // Parameters:
    //     AWLEN_param - The value to set onto wire <AWLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLEN( logic [3:0] AWLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLEN = AWLEN_param;
        else
            m_AWLEN <= AWLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWLEN_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWLEN_param - The value to set onto wire <AWLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLEN_index1( int _this_dot_1, logic  AWLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLEN[_this_dot_1] = AWLEN_param;
        else
            m_AWLEN[_this_dot_1] <= AWLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWLEN
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWLEN>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWLEN>.
    //
    function automatic logic [3:0]  get_AWLEN(  );
        return AWLEN;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWLEN_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWLEN>.
    //
    function automatic logic   get_AWLEN_index1( int _this_dot_1 );
        return AWLEN[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWSIZE
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWSIZE>.
    //
    // Parameters:
    //     AWSIZE_param - The value to set onto wire <AWSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWSIZE( logic [2:0] AWSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWSIZE = AWSIZE_param;
        else
            m_AWSIZE <= AWSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWSIZE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWSIZE_param - The value to set onto wire <AWSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWSIZE_index1( int _this_dot_1, logic  AWSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWSIZE[_this_dot_1] = AWSIZE_param;
        else
            m_AWSIZE[_this_dot_1] <= AWSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWSIZE
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWSIZE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWSIZE>.
    //
    function automatic logic [2:0]  get_AWSIZE(  );
        return AWSIZE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWSIZE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWSIZE>.
    //
    function automatic logic   get_AWSIZE_index1( int _this_dot_1 );
        return AWSIZE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWBURST
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWBURST>.
    //
    // Parameters:
    //     AWBURST_param - The value to set onto wire <AWBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWBURST( logic [1:0] AWBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWBURST = AWBURST_param;
        else
            m_AWBURST <= AWBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWBURST_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWBURST_param - The value to set onto wire <AWBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWBURST_index1( int _this_dot_1, logic  AWBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWBURST[_this_dot_1] = AWBURST_param;
        else
            m_AWBURST[_this_dot_1] <= AWBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWBURST
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWBURST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWBURST>.
    //
    function automatic logic [1:0]  get_AWBURST(  );
        return AWBURST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWBURST_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWBURST>.
    //
    function automatic logic   get_AWBURST_index1( int _this_dot_1 );
        return AWBURST[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWLOCK
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWLOCK>.
    //
    // Parameters:
    //     AWLOCK_param - The value to set onto wire <AWLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLOCK( logic [1:0] AWLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLOCK = AWLOCK_param;
        else
            m_AWLOCK <= AWLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWLOCK_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWLOCK_param - The value to set onto wire <AWLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLOCK_index1( int _this_dot_1, logic  AWLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLOCK[_this_dot_1] = AWLOCK_param;
        else
            m_AWLOCK[_this_dot_1] <= AWLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWLOCK
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWLOCK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWLOCK>.
    //
    function automatic logic [1:0]  get_AWLOCK(  );
        return AWLOCK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWLOCK_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWLOCK>.
    //
    function automatic logic   get_AWLOCK_index1( int _this_dot_1 );
        return AWLOCK[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWCACHE
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWCACHE>.
    //
    // Parameters:
    //     AWCACHE_param - The value to set onto wire <AWCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWCACHE( logic [3:0] AWCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWCACHE = AWCACHE_param;
        else
            m_AWCACHE <= AWCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWCACHE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWCACHE_param - The value to set onto wire <AWCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWCACHE_index1( int _this_dot_1, logic  AWCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWCACHE[_this_dot_1] = AWCACHE_param;
        else
            m_AWCACHE[_this_dot_1] <= AWCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWCACHE
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWCACHE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWCACHE>.
    //
    function automatic logic [3:0]  get_AWCACHE(  );
        return AWCACHE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWCACHE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWCACHE>.
    //
    function automatic logic   get_AWCACHE_index1( int _this_dot_1 );
        return AWCACHE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWPROT
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWPROT>.
    //
    // Parameters:
    //     AWPROT_param - The value to set onto wire <AWPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWPROT( logic [2:0] AWPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWPROT = AWPROT_param;
        else
            m_AWPROT <= AWPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWPROT_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWPROT_param - The value to set onto wire <AWPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWPROT_index1( int _this_dot_1, logic  AWPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWPROT[_this_dot_1] = AWPROT_param;
        else
            m_AWPROT[_this_dot_1] <= AWPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWPROT
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWPROT>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWPROT>.
    //
    function automatic logic [2:0]  get_AWPROT(  );
        return AWPROT;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWPROT_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWPROT>.
    //
    function automatic logic   get_AWPROT_index1( int _this_dot_1 );
        return AWPROT[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWID
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWID>.
    //
    // Parameters:
    //     AWID_param - The value to set onto wire <AWID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWID( logic [((AXI_ID_WIDTH) - 1):0]  AWID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWID = AWID_param;
        else
            m_AWID <= AWID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWID_param - The value to set onto wire <AWID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWID_index1( int _this_dot_1, logic  AWID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWID[_this_dot_1] = AWID_param;
        else
            m_AWID[_this_dot_1] <= AWID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWID
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_AWID(  );
        return AWID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWID>.
    //
    function automatic logic   get_AWID_index1( int _this_dot_1 );
        return AWID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWREADY>.
    //
    // Parameters:
    //     AWREADY_param - The value to set onto wire <AWREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWREADY( logic AWREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWREADY = AWREADY_param;
        else
            m_AWREADY <= AWREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWREADY>.
    //
    function automatic logic get_AWREADY(  );
        return AWREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWUSER>.
    //
    // Parameters:
    //     AWUSER_param - The value to set onto wire <AWUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWUSER( logic [7:0] AWUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWUSER = AWUSER_param;
        else
            m_AWUSER <= AWUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWUSER_param - The value to set onto wire <AWUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWUSER_index1( int _this_dot_1, logic  AWUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWUSER[_this_dot_1] = AWUSER_param;
        else
            m_AWUSER[_this_dot_1] <= AWUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWUSER>.
    //
    function automatic logic [7:0]  get_AWUSER(  );
        return AWUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWUSER>.
    //
    function automatic logic   get_AWUSER_index1( int _this_dot_1 );
        return AWUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARVALID>.
    //
    // Parameters:
    //     ARVALID_param - The value to set onto wire <ARVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARVALID( logic ARVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARVALID = ARVALID_param;
        else
            m_ARVALID <= ARVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARVALID>.
    //
    function automatic logic get_ARVALID(  );
        return ARVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARADDR
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARADDR>.
    //
    // Parameters:
    //     ARADDR_param - The value to set onto wire <ARADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARADDR( logic [((AXI_ADDRESS_WIDTH) - 1):0]  ARADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARADDR = ARADDR_param;
        else
            m_ARADDR <= ARADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARADDR_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARADDR_param - The value to set onto wire <ARADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARADDR_index1( int _this_dot_1, logic  ARADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARADDR[_this_dot_1] = ARADDR_param;
        else
            m_ARADDR[_this_dot_1] <= ARADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARADDR
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARADDR>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARADDR>.
    //
    function automatic logic [((AXI_ADDRESS_WIDTH) - 1):0]   get_ARADDR(  );
        return ARADDR;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARADDR_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARADDR>.
    //
    function automatic logic   get_ARADDR_index1( int _this_dot_1 );
        return ARADDR[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARLEN
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARLEN>.
    //
    // Parameters:
    //     ARLEN_param - The value to set onto wire <ARLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLEN( logic [3:0] ARLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLEN = ARLEN_param;
        else
            m_ARLEN <= ARLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARLEN_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARLEN_param - The value to set onto wire <ARLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLEN_index1( int _this_dot_1, logic  ARLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLEN[_this_dot_1] = ARLEN_param;
        else
            m_ARLEN[_this_dot_1] <= ARLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARLEN
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARLEN>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARLEN>.
    //
    function automatic logic [3:0]  get_ARLEN(  );
        return ARLEN;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARLEN_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARLEN>.
    //
    function automatic logic   get_ARLEN_index1( int _this_dot_1 );
        return ARLEN[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARSIZE
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARSIZE>.
    //
    // Parameters:
    //     ARSIZE_param - The value to set onto wire <ARSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARSIZE( logic [2:0] ARSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARSIZE = ARSIZE_param;
        else
            m_ARSIZE <= ARSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARSIZE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARSIZE_param - The value to set onto wire <ARSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARSIZE_index1( int _this_dot_1, logic  ARSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARSIZE[_this_dot_1] = ARSIZE_param;
        else
            m_ARSIZE[_this_dot_1] <= ARSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARSIZE
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARSIZE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARSIZE>.
    //
    function automatic logic [2:0]  get_ARSIZE(  );
        return ARSIZE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARSIZE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARSIZE>.
    //
    function automatic logic   get_ARSIZE_index1( int _this_dot_1 );
        return ARSIZE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARBURST
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARBURST>.
    //
    // Parameters:
    //     ARBURST_param - The value to set onto wire <ARBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARBURST( logic [1:0] ARBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARBURST = ARBURST_param;
        else
            m_ARBURST <= ARBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARBURST_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARBURST_param - The value to set onto wire <ARBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARBURST_index1( int _this_dot_1, logic  ARBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARBURST[_this_dot_1] = ARBURST_param;
        else
            m_ARBURST[_this_dot_1] <= ARBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARBURST
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARBURST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARBURST>.
    //
    function automatic logic [1:0]  get_ARBURST(  );
        return ARBURST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARBURST_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARBURST>.
    //
    function automatic logic   get_ARBURST_index1( int _this_dot_1 );
        return ARBURST[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARLOCK
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARLOCK>.
    //
    // Parameters:
    //     ARLOCK_param - The value to set onto wire <ARLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLOCK( logic [1:0] ARLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLOCK = ARLOCK_param;
        else
            m_ARLOCK <= ARLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARLOCK_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARLOCK_param - The value to set onto wire <ARLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLOCK_index1( int _this_dot_1, logic  ARLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLOCK[_this_dot_1] = ARLOCK_param;
        else
            m_ARLOCK[_this_dot_1] <= ARLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARLOCK
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARLOCK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARLOCK>.
    //
    function automatic logic [1:0]  get_ARLOCK(  );
        return ARLOCK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARLOCK_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARLOCK>.
    //
    function automatic logic   get_ARLOCK_index1( int _this_dot_1 );
        return ARLOCK[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARCACHE
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARCACHE>.
    //
    // Parameters:
    //     ARCACHE_param - The value to set onto wire <ARCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARCACHE( logic [3:0] ARCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARCACHE = ARCACHE_param;
        else
            m_ARCACHE <= ARCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARCACHE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARCACHE_param - The value to set onto wire <ARCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARCACHE_index1( int _this_dot_1, logic  ARCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARCACHE[_this_dot_1] = ARCACHE_param;
        else
            m_ARCACHE[_this_dot_1] <= ARCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARCACHE
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARCACHE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARCACHE>.
    //
    function automatic logic [3:0]  get_ARCACHE(  );
        return ARCACHE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARCACHE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARCACHE>.
    //
    function automatic logic   get_ARCACHE_index1( int _this_dot_1 );
        return ARCACHE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARPROT
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARPROT>.
    //
    // Parameters:
    //     ARPROT_param - The value to set onto wire <ARPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARPROT( logic [2:0] ARPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARPROT = ARPROT_param;
        else
            m_ARPROT <= ARPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARPROT_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARPROT_param - The value to set onto wire <ARPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARPROT_index1( int _this_dot_1, logic  ARPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARPROT[_this_dot_1] = ARPROT_param;
        else
            m_ARPROT[_this_dot_1] <= ARPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARPROT
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARPROT>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARPROT>.
    //
    function automatic logic [2:0]  get_ARPROT(  );
        return ARPROT;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARPROT_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARPROT>.
    //
    function automatic logic   get_ARPROT_index1( int _this_dot_1 );
        return ARPROT[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARID
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARID>.
    //
    // Parameters:
    //     ARID_param - The value to set onto wire <ARID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARID( logic [((AXI_ID_WIDTH) - 1):0]  ARID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARID = ARID_param;
        else
            m_ARID <= ARID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARID_param - The value to set onto wire <ARID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARID_index1( int _this_dot_1, logic  ARID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARID[_this_dot_1] = ARID_param;
        else
            m_ARID[_this_dot_1] <= ARID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARID
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_ARID(  );
        return ARID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARID>.
    //
    function automatic logic   get_ARID_index1( int _this_dot_1 );
        return ARID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARREADY>.
    //
    // Parameters:
    //     ARREADY_param - The value to set onto wire <ARREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARREADY( logic ARREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARREADY = ARREADY_param;
        else
            m_ARREADY <= ARREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARREADY>.
    //
    function automatic logic get_ARREADY(  );
        return ARREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARUSER>.
    //
    // Parameters:
    //     ARUSER_param - The value to set onto wire <ARUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARUSER( logic [7:0] ARUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARUSER = ARUSER_param;
        else
            m_ARUSER <= ARUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARUSER_param - The value to set onto wire <ARUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARUSER_index1( int _this_dot_1, logic  ARUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARUSER[_this_dot_1] = ARUSER_param;
        else
            m_ARUSER[_this_dot_1] <= ARUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARUSER>.
    //
    function automatic logic [7:0]  get_ARUSER(  );
        return ARUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARUSER>.
    //
    function automatic logic   get_ARUSER_index1( int _this_dot_1 );
        return ARUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <RVALID>.
    //
    // Parameters:
    //     RVALID_param - The value to set onto wire <RVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RVALID( logic RVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RVALID = RVALID_param;
        else
            m_RVALID <= RVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <RVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RVALID>.
    //
    function automatic logic get_RVALID(  );
        return RVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RLAST
    //-------------------------------------------------------------------------
    //     Set the value of wire <RLAST>.
    //
    // Parameters:
    //     RLAST_param - The value to set onto wire <RLAST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RLAST( logic RLAST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RLAST = RLAST_param;
        else
            m_RLAST <= RLAST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RLAST
    //-------------------------------------------------------------------------
    //     Get the value of wire <RLAST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RLAST>.
    //
    function automatic logic get_RLAST(  );
        return RLAST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RDATA
    //-------------------------------------------------------------------------
    //     Set the value of wire <RDATA>.
    //
    // Parameters:
    //     RDATA_param - The value to set onto wire <RDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RDATA( logic [((AXI_RDATA_WIDTH) - 1):0]  RDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RDATA = RDATA_param;
        else
            m_RDATA <= RDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RDATA_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RDATA_param - The value to set onto wire <RDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RDATA_index1( int _this_dot_1, logic  RDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RDATA[_this_dot_1] = RDATA_param;
        else
            m_RDATA[_this_dot_1] <= RDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RDATA
    //-------------------------------------------------------------------------
    //     Get the value of wire <RDATA>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RDATA>.
    //
    function automatic logic [((AXI_RDATA_WIDTH) - 1):0]   get_RDATA(  );
        return RDATA;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RDATA_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RDATA>.
    //
    function automatic logic   get_RDATA_index1( int _this_dot_1 );
        return RDATA[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RRESP
    //-------------------------------------------------------------------------
    //     Set the value of wire <RRESP>.
    //
    // Parameters:
    //     RRESP_param - The value to set onto wire <RRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RRESP( logic [1:0] RRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RRESP = RRESP_param;
        else
            m_RRESP <= RRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RRESP_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RRESP_param - The value to set onto wire <RRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RRESP_index1( int _this_dot_1, logic  RRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RRESP[_this_dot_1] = RRESP_param;
        else
            m_RRESP[_this_dot_1] <= RRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RRESP
    //-------------------------------------------------------------------------
    //     Get the value of wire <RRESP>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RRESP>.
    //
    function automatic logic [1:0]  get_RRESP(  );
        return RRESP;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RRESP_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RRESP>.
    //
    function automatic logic   get_RRESP_index1( int _this_dot_1 );
        return RRESP[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RID
    //-------------------------------------------------------------------------
    //     Set the value of wire <RID>.
    //
    // Parameters:
    //     RID_param - The value to set onto wire <RID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RID( logic [((AXI_ID_WIDTH) - 1):0]  RID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RID = RID_param;
        else
            m_RID <= RID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RID_param - The value to set onto wire <RID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RID_index1( int _this_dot_1, logic  RID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RID[_this_dot_1] = RID_param;
        else
            m_RID[_this_dot_1] <= RID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RID
    //-------------------------------------------------------------------------
    //     Get the value of wire <RID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_RID(  );
        return RID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RID>.
    //
    function automatic logic   get_RID_index1( int _this_dot_1 );
        return RID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <RREADY>.
    //
    // Parameters:
    //     RREADY_param - The value to set onto wire <RREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RREADY( logic RREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RREADY = RREADY_param;
        else
            m_RREADY <= RREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <RREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RREADY>.
    //
    function automatic logic get_RREADY(  );
        return RREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <RUSER>.
    //
    // Parameters:
    //     RUSER_param - The value to set onto wire <RUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RUSER( logic [7:0] RUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RUSER = RUSER_param;
        else
            m_RUSER <= RUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RUSER_param - The value to set onto wire <RUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RUSER_index1( int _this_dot_1, logic  RUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RUSER[_this_dot_1] = RUSER_param;
        else
            m_RUSER[_this_dot_1] <= RUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <RUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RUSER>.
    //
    function automatic logic [7:0]  get_RUSER(  );
        return RUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RUSER>.
    //
    function automatic logic   get_RUSER_index1( int _this_dot_1 );
        return RUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <WVALID>.
    //
    // Parameters:
    //     WVALID_param - The value to set onto wire <WVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WVALID( logic WVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WVALID = WVALID_param;
        else
            m_WVALID <= WVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <WVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WVALID>.
    //
    function automatic logic get_WVALID(  );
        return WVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WLAST
    //-------------------------------------------------------------------------
    //     Set the value of wire <WLAST>.
    //
    // Parameters:
    //     WLAST_param - The value to set onto wire <WLAST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WLAST( logic WLAST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WLAST = WLAST_param;
        else
            m_WLAST <= WLAST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WLAST
    //-------------------------------------------------------------------------
    //     Get the value of wire <WLAST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WLAST>.
    //
    function automatic logic get_WLAST(  );
        return WLAST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WDATA
    //-------------------------------------------------------------------------
    //     Set the value of wire <WDATA>.
    //
    // Parameters:
    //     WDATA_param - The value to set onto wire <WDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WDATA( logic [((AXI_WDATA_WIDTH) - 1):0]  WDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WDATA = WDATA_param;
        else
            m_WDATA <= WDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WDATA_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WDATA_param - The value to set onto wire <WDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WDATA_index1( int _this_dot_1, logic  WDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WDATA[_this_dot_1] = WDATA_param;
        else
            m_WDATA[_this_dot_1] <= WDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WDATA
    //-------------------------------------------------------------------------
    //     Get the value of wire <WDATA>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WDATA>.
    //
    function automatic logic [((AXI_WDATA_WIDTH) - 1):0]   get_WDATA(  );
        return WDATA;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WDATA_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WDATA>.
    //
    function automatic logic   get_WDATA_index1( int _this_dot_1 );
        return WDATA[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WSTRB
    //-------------------------------------------------------------------------
    //     Set the value of wire <WSTRB>.
    //
    // Parameters:
    //     WSTRB_param - The value to set onto wire <WSTRB>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WSTRB( logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  WSTRB_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WSTRB = WSTRB_param;
        else
            m_WSTRB <= WSTRB_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WSTRB_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WSTRB>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WSTRB_param - The value to set onto wire <WSTRB>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WSTRB_index1( int _this_dot_1, logic  WSTRB_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WSTRB[_this_dot_1] = WSTRB_param;
        else
            m_WSTRB[_this_dot_1] <= WSTRB_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WSTRB
    //-------------------------------------------------------------------------
    //     Get the value of wire <WSTRB>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WSTRB>.
    //
    function automatic logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]   get_WSTRB(  );
        return WSTRB;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WSTRB_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WSTRB>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WSTRB>.
    //
    function automatic logic   get_WSTRB_index1( int _this_dot_1 );
        return WSTRB[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WID
    //-------------------------------------------------------------------------
    //     Set the value of wire <WID>.
    //
    // Parameters:
    //     WID_param - The value to set onto wire <WID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WID( logic [((AXI_ID_WIDTH) - 1):0]  WID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WID = WID_param;
        else
            m_WID <= WID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WID_param - The value to set onto wire <WID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WID_index1( int _this_dot_1, logic  WID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WID[_this_dot_1] = WID_param;
        else
            m_WID[_this_dot_1] <= WID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WID
    //-------------------------------------------------------------------------
    //     Get the value of wire <WID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_WID(  );
        return WID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WID>.
    //
    function automatic logic   get_WID_index1( int _this_dot_1 );
        return WID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <WREADY>.
    //
    // Parameters:
    //     WREADY_param - The value to set onto wire <WREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WREADY( logic WREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WREADY = WREADY_param;
        else
            m_WREADY <= WREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <WREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WREADY>.
    //
    function automatic logic get_WREADY(  );
        return WREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <WUSER>.
    //
    // Parameters:
    //     WUSER_param - The value to set onto wire <WUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WUSER( logic [7:0] WUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WUSER = WUSER_param;
        else
            m_WUSER <= WUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WUSER_param - The value to set onto wire <WUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WUSER_index1( int _this_dot_1, logic  WUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WUSER[_this_dot_1] = WUSER_param;
        else
            m_WUSER[_this_dot_1] <= WUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <WUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WUSER>.
    //
    function automatic logic [7:0]  get_WUSER(  );
        return WUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WUSER>.
    //
    function automatic logic   get_WUSER_index1( int _this_dot_1 );
        return WUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <BVALID>.
    //
    // Parameters:
    //     BVALID_param - The value to set onto wire <BVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BVALID( logic BVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BVALID = BVALID_param;
        else
            m_BVALID <= BVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <BVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BVALID>.
    //
    function automatic logic get_BVALID(  );
        return BVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BRESP
    //-------------------------------------------------------------------------
    //     Set the value of wire <BRESP>.
    //
    // Parameters:
    //     BRESP_param - The value to set onto wire <BRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BRESP( logic [1:0] BRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BRESP = BRESP_param;
        else
            m_BRESP <= BRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BRESP_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BRESP_param - The value to set onto wire <BRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BRESP_index1( int _this_dot_1, logic  BRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BRESP[_this_dot_1] = BRESP_param;
        else
            m_BRESP[_this_dot_1] <= BRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BRESP
    //-------------------------------------------------------------------------
    //     Get the value of wire <BRESP>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BRESP>.
    //
    function automatic logic [1:0]  get_BRESP(  );
        return BRESP;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BRESP_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BRESP>.
    //
    function automatic logic   get_BRESP_index1( int _this_dot_1 );
        return BRESP[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BID
    //-------------------------------------------------------------------------
    //     Set the value of wire <BID>.
    //
    // Parameters:
    //     BID_param - The value to set onto wire <BID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BID( logic [((AXI_ID_WIDTH) - 1):0]  BID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BID = BID_param;
        else
            m_BID <= BID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BID_param - The value to set onto wire <BID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BID_index1( int _this_dot_1, logic  BID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BID[_this_dot_1] = BID_param;
        else
            m_BID[_this_dot_1] <= BID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BID
    //-------------------------------------------------------------------------
    //     Get the value of wire <BID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_BID(  );
        return BID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BID>.
    //
    function automatic logic   get_BID_index1( int _this_dot_1 );
        return BID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <BREADY>.
    //
    // Parameters:
    //     BREADY_param - The value to set onto wire <BREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BREADY( logic BREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BREADY = BREADY_param;
        else
            m_BREADY <= BREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <BREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BREADY>.
    //
    function automatic logic get_BREADY(  );
        return BREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <BUSER>.
    //
    // Parameters:
    //     BUSER_param - The value to set onto wire <BUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BUSER( logic [7:0] BUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BUSER = BUSER_param;
        else
            m_BUSER <= BUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BUSER_param - The value to set onto wire <BUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BUSER_index1( int _this_dot_1, logic  BUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BUSER[_this_dot_1] = BUSER_param;
        else
            m_BUSER[_this_dot_1] <= BUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <BUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BUSER>.
    //
    function automatic logic [7:0]  get_BUSER(  );
        return BUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BUSER>.
    //
    function automatic logic   get_BUSER_index1( int _this_dot_1 );
        return BUSER[_this_dot_1];
    endfunction

    //-------------------------------------------------------------------------
    // Tasks to wait for a change to a global variable with read access
    //-------------------------------------------------------------------------


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_write_ctrl_to_data_mintime
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_write_ctrl_to_data_mintime>.
    //
    task automatic wait_for_config_write_ctrl_to_data_mintime(  );
        begin
            @( config_write_ctrl_to_data_mintime );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_master_write_delay
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_master_write_delay>.
    //
    task automatic wait_for_config_master_write_delay(  );
        begin
            @( config_master_write_delay );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_all_assertions
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_all_assertions>.
    //
    task automatic wait_for_config_enable_all_assertions(  );
        begin
            @( config_enable_all_assertions );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_assertion
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_assertion>.
    //
    task automatic wait_for_config_enable_assertion(  );
        begin
            @( config_enable_assertion );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_assertion_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_enable_assertion_index1( input int _this_dot_1 );
        begin
            @( config_enable_assertion[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_start_addr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_start_addr>.
    //
    task automatic wait_for_config_slave_start_addr(  );
        begin
            @( config_slave_start_addr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_start_addr_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_slave_start_addr_index1( input int _this_dot_1 );
        begin
            @( config_slave_start_addr[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_end_addr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_end_addr>.
    //
    task automatic wait_for_config_slave_end_addr(  );
        begin
            @( config_slave_end_addr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_end_addr_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_slave_end_addr_index1( input int _this_dot_1 );
        begin
            @( config_slave_end_addr[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_support_exclusive_access
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_support_exclusive_access>.
    //
    task automatic wait_for_config_support_exclusive_access(  );
        begin
            @( config_support_exclusive_access );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_read_data_reordering_depth
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_read_data_reordering_depth>.
    //
    task automatic wait_for_config_read_data_reordering_depth(  );
        begin
            @( config_read_data_reordering_depth );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_transaction_time_factor
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_transaction_time_factor>.
    //
    task automatic wait_for_config_max_transaction_time_factor(  );
        begin
            @( config_max_transaction_time_factor );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_timeout_max_data_transfer
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_timeout_max_data_transfer>.
    //
    task automatic wait_for_config_timeout_max_data_transfer(  );
        begin
            @( config_timeout_max_data_transfer );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_burst_timeout_factor
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_burst_timeout_factor>.
    //
    task automatic wait_for_config_burst_timeout_factor(  );
        begin
            @( config_burst_timeout_factor );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_AWVALID_assertion_to_AWREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    task automatic wait_for_config_max_latency_AWVALID_assertion_to_AWREADY(  );
        begin
            @( config_max_latency_AWVALID_assertion_to_AWREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_ARVALID_assertion_to_ARREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    task automatic wait_for_config_max_latency_ARVALID_assertion_to_ARREADY(  );
        begin
            @( config_max_latency_ARVALID_assertion_to_ARREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_RVALID_assertion_to_RREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_RVALID_assertion_to_RREADY>.
    //
    task automatic wait_for_config_max_latency_RVALID_assertion_to_RREADY(  );
        begin
            @( config_max_latency_RVALID_assertion_to_RREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_BVALID_assertion_to_BREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_BVALID_assertion_to_BREADY>.
    //
    task automatic wait_for_config_max_latency_BVALID_assertion_to_BREADY(  );
        begin
            @( config_max_latency_BVALID_assertion_to_BREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_WVALID_assertion_to_WREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_WVALID_assertion_to_WREADY>.
    //
    task automatic wait_for_config_max_latency_WVALID_assertion_to_WREADY(  );
        begin
            @( config_max_latency_WVALID_assertion_to_WREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_master_error_position
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_master_error_position>.
    //
    task automatic wait_for_config_master_error_position(  );
        begin
            @( config_master_error_position );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_setup_time
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_setup_time>.
    //
    task automatic wait_for_config_setup_time(  );
        begin
            @( config_setup_time );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_hold_time
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_hold_time>.
    //
    task automatic wait_for_config_hold_time(  );
        begin
            @( config_hold_time );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_wr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_wr>.
    //
    task automatic wait_for_config_max_outstanding_wr(  );
        begin
            @( config_max_outstanding_wr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_rd
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_rd>.
    //
    task automatic wait_for_config_max_outstanding_rd(  );
        begin
            @( config_max_outstanding_rd );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_rw
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_rw>.
    //
    task automatic wait_for_config_max_outstanding_rw(  );
        begin
            @( config_max_outstanding_rw );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_is_issuing
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_is_issuing>.
    //
    task automatic wait_for_config_is_issuing(  );
        begin
            @( config_is_issuing );
        end
    endtask


    //-------------------------------------------------------------------------
    // Functions to set global variables with write access
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- set_config_write_ctrl_to_data_mintime
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_write_ctrl_to_data_mintime>.
    //
    // Parameters:
    //     config_write_ctrl_to_data_mintime_param - The value to assign to variable <config_write_ctrl_to_data_mintime>.
    //
    function automatic void set_config_write_ctrl_to_data_mintime( int unsigned config_write_ctrl_to_data_mintime_param );
        config_write_ctrl_to_data_mintime = config_write_ctrl_to_data_mintime_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_master_write_delay
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_master_write_delay>.
    //
    // Parameters:
    //     config_master_write_delay_param - The value to assign to variable <config_master_write_delay>.
    //
    function automatic void set_config_master_write_delay( bit config_master_write_delay_param );
        config_master_write_delay = config_master_write_delay_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_all_assertions
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_enable_all_assertions>.
    //
    // Parameters:
    //     config_enable_all_assertions_param - The value to assign to variable <config_enable_all_assertions>.
    //
    function automatic void set_config_enable_all_assertions( bit config_enable_all_assertions_param );
        config_enable_all_assertions = config_enable_all_assertions_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_assertion
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_enable_assertion>.
    //
    // Parameters:
    //     config_enable_assertion_param - The value to assign to variable <config_enable_assertion>.
    //
    function automatic void set_config_enable_assertion( bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
        config_enable_assertion = config_enable_assertion_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_assertion_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_enable_assertion_param - The value to assign to variable <config_enable_assertion>.
    //
    function automatic void set_config_enable_assertion_index1( int _this_dot_1, bit  config_enable_assertion_param );
        config_enable_assertion[_this_dot_1] = config_enable_assertion_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_start_addr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_slave_start_addr>.
    //
    // Parameters:
    //     config_slave_start_addr_param - The value to assign to variable <config_slave_start_addr>.
    //
    function automatic void set_config_slave_start_addr( bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param );
        config_slave_start_addr = config_slave_start_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_start_addr_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_slave_start_addr_param - The value to assign to variable <config_slave_start_addr>.
    //
    function automatic void set_config_slave_start_addr_index1( int _this_dot_1, bit  config_slave_start_addr_param );
        config_slave_start_addr[_this_dot_1] = config_slave_start_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_end_addr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_slave_end_addr>.
    //
    // Parameters:
    //     config_slave_end_addr_param - The value to assign to variable <config_slave_end_addr>.
    //
    function automatic void set_config_slave_end_addr( bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param );
        config_slave_end_addr = config_slave_end_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_end_addr_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_slave_end_addr_param - The value to assign to variable <config_slave_end_addr>.
    //
    function automatic void set_config_slave_end_addr_index1( int _this_dot_1, bit  config_slave_end_addr_param );
        config_slave_end_addr[_this_dot_1] = config_slave_end_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_support_exclusive_access
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_support_exclusive_access>.
    //
    // Parameters:
    //     config_support_exclusive_access_param - The value to assign to variable <config_support_exclusive_access>.
    //
    function automatic void set_config_support_exclusive_access( bit config_support_exclusive_access_param );
        config_support_exclusive_access = config_support_exclusive_access_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_read_data_reordering_depth
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_read_data_reordering_depth>.
    //
    // Parameters:
    //     config_read_data_reordering_depth_param - The value to assign to variable <config_read_data_reordering_depth>.
    //
    function automatic void set_config_read_data_reordering_depth( int unsigned config_read_data_reordering_depth_param );
        config_read_data_reordering_depth = config_read_data_reordering_depth_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_transaction_time_factor
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_transaction_time_factor>.
    //
    // Parameters:
    //     config_max_transaction_time_factor_param - The value to assign to variable <config_max_transaction_time_factor>.
    //
    function automatic void set_config_max_transaction_time_factor( int unsigned config_max_transaction_time_factor_param );
        config_max_transaction_time_factor = config_max_transaction_time_factor_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_timeout_max_data_transfer
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_timeout_max_data_transfer>.
    //
    // Parameters:
    //     config_timeout_max_data_transfer_param - The value to assign to variable <config_timeout_max_data_transfer>.
    //
    function automatic void set_config_timeout_max_data_transfer( int config_timeout_max_data_transfer_param );
        config_timeout_max_data_transfer = config_timeout_max_data_transfer_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_burst_timeout_factor
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_burst_timeout_factor>.
    //
    // Parameters:
    //     config_burst_timeout_factor_param - The value to assign to variable <config_burst_timeout_factor>.
    //
    function automatic void set_config_burst_timeout_factor( int unsigned config_burst_timeout_factor_param );
        config_burst_timeout_factor = config_burst_timeout_factor_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_AWVALID_assertion_to_AWREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    // Parameters:
    //     config_max_latency_AWVALID_assertion_to_AWREADY_param - The value to assign to variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    function automatic void set_config_max_latency_AWVALID_assertion_to_AWREADY( int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
        config_max_latency_AWVALID_assertion_to_AWREADY = config_max_latency_AWVALID_assertion_to_AWREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_ARVALID_assertion_to_ARREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    // Parameters:
    //     config_max_latency_ARVALID_assertion_to_ARREADY_param - The value to assign to variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    function automatic void set_config_max_latency_ARVALID_assertion_to_ARREADY( int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
        config_max_latency_ARVALID_assertion_to_ARREADY = config_max_latency_ARVALID_assertion_to_ARREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_RVALID_assertion_to_RREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    // Parameters:
    //     config_max_latency_RVALID_assertion_to_RREADY_param - The value to assign to variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    function automatic void set_config_max_latency_RVALID_assertion_to_RREADY( int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
        config_max_latency_RVALID_assertion_to_RREADY = config_max_latency_RVALID_assertion_to_RREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_BVALID_assertion_to_BREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    // Parameters:
    //     config_max_latency_BVALID_assertion_to_BREADY_param - The value to assign to variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    function automatic void set_config_max_latency_BVALID_assertion_to_BREADY( int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
        config_max_latency_BVALID_assertion_to_BREADY = config_max_latency_BVALID_assertion_to_BREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_WVALID_assertion_to_WREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    // Parameters:
    //     config_max_latency_WVALID_assertion_to_WREADY_param - The value to assign to variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    function automatic void set_config_max_latency_WVALID_assertion_to_WREADY( int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
        config_max_latency_WVALID_assertion_to_WREADY = config_max_latency_WVALID_assertion_to_WREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_master_error_position
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_master_error_position>.
    //
    // Parameters:
    //     config_master_error_position_param - The value to assign to variable <config_master_error_position>.
    //
    function automatic void set_config_master_error_position( axi_error_e config_master_error_position_param );
        config_master_error_position = config_master_error_position_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_setup_time
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_setup_time>.
    //
    // Parameters:
    //     config_setup_time_param - The value to assign to variable <config_setup_time>.
    //
    function automatic void set_config_setup_time( int config_setup_time_param );
        config_setup_time = config_setup_time_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_hold_time
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_hold_time>.
    //
    // Parameters:
    //     config_hold_time_param - The value to assign to variable <config_hold_time>.
    //
    function automatic void set_config_hold_time( int config_hold_time_param );
        config_hold_time = config_hold_time_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_wr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_wr>.
    //
    // Parameters:
    //     config_max_outstanding_wr_param - The value to assign to variable <config_max_outstanding_wr>.
    //
    function automatic void set_config_max_outstanding_wr( int config_max_outstanding_wr_param );
        config_max_outstanding_wr = config_max_outstanding_wr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_rd
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_rd>.
    //
    // Parameters:
    //     config_max_outstanding_rd_param - The value to assign to variable <config_max_outstanding_rd>.
    //
    function automatic void set_config_max_outstanding_rd( int config_max_outstanding_rd_param );
        config_max_outstanding_rd = config_max_outstanding_rd_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_rw
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_rw>.
    //
    // Parameters:
    //     config_max_outstanding_rw_param - The value to assign to variable <config_max_outstanding_rw>.
    //
    function automatic void set_config_max_outstanding_rw( int config_max_outstanding_rw_param );
        config_max_outstanding_rw = config_max_outstanding_rw_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_is_issuing
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_is_issuing>.
    //
    // Parameters:
    //     config_is_issuing_param - The value to assign to variable <config_is_issuing>.
    //
    function automatic void set_config_is_issuing( bit config_is_issuing_param );
        config_is_issuing = config_is_issuing_param;
    endfunction


    //-------------------------------------------------------------------------
    // Functions to get global variables with read access
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- get_config_write_ctrl_to_data_mintime
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_write_ctrl_to_data_mintime>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_write_ctrl_to_data_mintime>.
    //
    function automatic int unsigned get_config_write_ctrl_to_data_mintime(  );
        return config_write_ctrl_to_data_mintime;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_master_write_delay
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_master_write_delay>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_master_write_delay>.
    //
    function automatic bit get_config_master_write_delay(  );
        axi_get_deprecated_config_master_write_delay_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_master_write_delay;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_all_assertions
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_enable_all_assertions>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_enable_all_assertions>.
    //
    function automatic bit get_config_enable_all_assertions(  );
        return config_enable_all_assertions;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_assertion
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_enable_assertion>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_enable_assertion>.
    //
    function automatic bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]   get_config_enable_assertion(  );
        return config_enable_assertion;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_assertion_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_enable_assertion>.
    //
    function automatic bit   get_config_enable_assertion_index1( int _this_dot_1 );
        return config_enable_assertion[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_start_addr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_slave_start_addr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_slave_start_addr>.
    //
    function automatic bit [((AXI_ADDRESS_WIDTH) - 1):0]   get_config_slave_start_addr(  );
        axi_get_deprecated_config_slave_start_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_start_addr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_start_addr_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_slave_start_addr>.
    //
    function automatic bit   get_config_slave_start_addr_index1( int _this_dot_1 );
        axi_get_deprecated_config_slave_start_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_start_addr[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_end_addr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_slave_end_addr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_slave_end_addr>.
    //
    function automatic bit [((AXI_ADDRESS_WIDTH) - 1):0]   get_config_slave_end_addr(  );
        axi_get_deprecated_config_slave_end_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_end_addr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_end_addr_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_slave_end_addr>.
    //
    function automatic bit   get_config_slave_end_addr_index1( int _this_dot_1 );
        axi_get_deprecated_config_slave_end_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_end_addr[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_support_exclusive_access
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_support_exclusive_access>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_support_exclusive_access>.
    //
    function automatic bit get_config_support_exclusive_access(  );
        return config_support_exclusive_access;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_read_data_reordering_depth
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_read_data_reordering_depth>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_read_data_reordering_depth>.
    //
    function automatic int unsigned get_config_read_data_reordering_depth(  );
        return config_read_data_reordering_depth;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_transaction_time_factor
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_transaction_time_factor>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_transaction_time_factor>.
    //
    function automatic int unsigned get_config_max_transaction_time_factor(  );
        return config_max_transaction_time_factor;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_timeout_max_data_transfer
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_timeout_max_data_transfer>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_timeout_max_data_transfer>.
    //
    function automatic int get_config_timeout_max_data_transfer(  );
        return config_timeout_max_data_transfer;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_burst_timeout_factor
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_burst_timeout_factor>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_burst_timeout_factor>.
    //
    function automatic int unsigned get_config_burst_timeout_factor(  );
        return config_burst_timeout_factor;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_AWVALID_assertion_to_AWREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    function automatic int unsigned get_config_max_latency_AWVALID_assertion_to_AWREADY(  );
        return config_max_latency_AWVALID_assertion_to_AWREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_ARVALID_assertion_to_ARREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    function automatic int unsigned get_config_max_latency_ARVALID_assertion_to_ARREADY(  );
        return config_max_latency_ARVALID_assertion_to_ARREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_RVALID_assertion_to_RREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    function automatic int unsigned get_config_max_latency_RVALID_assertion_to_RREADY(  );
        return config_max_latency_RVALID_assertion_to_RREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_BVALID_assertion_to_BREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    function automatic int unsigned get_config_max_latency_BVALID_assertion_to_BREADY(  );
        return config_max_latency_BVALID_assertion_to_BREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_WVALID_assertion_to_WREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    function automatic int unsigned get_config_max_latency_WVALID_assertion_to_WREADY(  );
        return config_max_latency_WVALID_assertion_to_WREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_master_error_position
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_master_error_position>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_master_error_position>.
    //
    function automatic axi_error_e get_config_master_error_position(  );
        axi_get_deprecated_config_master_error_position_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_master_error_position;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_setup_time
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_setup_time>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_setup_time>.
    //
    function automatic int get_config_setup_time(  );
        return config_setup_time;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_hold_time
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_hold_time>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_hold_time>.
    //
    function automatic int get_config_hold_time(  );
        return config_hold_time;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_wr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_wr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_wr>.
    //
    function automatic int get_config_max_outstanding_wr(  );
        return config_max_outstanding_wr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_rd
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_rd>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_rd>.
    //
    function automatic int get_config_max_outstanding_rd(  );
        return config_max_outstanding_rd;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_rw
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_rw>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_rw>.
    //
    function automatic int get_config_max_outstanding_rw(  );
        return config_max_outstanding_rw;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_is_issuing
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_is_issuing>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_is_issuing>.
    //
    function automatic bit get_config_is_issuing(  );
        return config_is_issuing;
    endfunction


    //-------------------------------------------------------------------------
    // Functions to set/get generic interface configuration
    //-------------------------------------------------------------------------

    function void set_interface
    (
        input int what = 0,
        input int arg1 = 0,
        input int arg2 = 0,
        input int arg3 = 0,
        input int arg4 = 0,
        input int arg5 = 0,
        input int arg6 = 0,
        input int arg7 = 0,
        input int arg8 = 0,
        input int arg9 = 0,
        input int arg10 = 0
    );
        axi_set_interface( what, arg1, arg2, arg3, arg4, arg5, arg6, arg7, arg8, arg9, arg10 );
    endfunction

    function int get_interface
    (
        input int what = 0,
        input int arg1 = 0,
        input int arg2 = 0,
        input int arg3 = 0,
        input int arg4 = 0,
        input int arg5 = 0,
        input int arg6 = 0,
        input int arg7 = 0,
        input int arg8 = 0,
        input int arg9 = 0
    );
        return axi_get_interface( what, arg1, arg2, arg3, arg4, arg5, arg6, arg7, arg8, arg9 );
    endfunction

    //-------------------------------------------------------------------------
    // Functions to get the hierarchic name of this interface
    //-------------------------------------------------------------------------
    function string get_full_name();
        return axi_get_full_name();
    endfunction

    //--------------------------------------------------------------------------
    //
    // Group:- Monitor Value Change on Variable
    //
    //--------------------------------------------------------------------------

    function automatic void axi_local_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( ref int unsigned config_write_ctrl_to_data_mintime_param );
        axi_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( _interface_ref, config_write_ctrl_to_data_mintime );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( config_write_ctrl_to_data_mintime );
            end
        end
    end

    function automatic void axi_local_set_config_master_write_delay_from_SystemVerilog( ref bit config_master_write_delay_param );
        axi_set_config_master_write_delay_from_SystemVerilog( _interface_ref, config_master_write_delay );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_master_write_delay_from_SystemVerilog( config_master_write_delay );
            end
        end
    end

    function automatic void axi_local_set_config_enable_all_assertions_from_SystemVerilog( ref bit config_enable_all_assertions_param );
        axi_set_config_enable_all_assertions_from_SystemVerilog( _interface_ref, config_enable_all_assertions );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_enable_all_assertions_from_SystemVerilog( config_enable_all_assertions );
            end
        end
    end

    function automatic void axi_local_set_config_enable_assertion_from_SystemVerilog( ref bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
        axi_set_config_enable_assertion_from_SystemVerilog( _interface_ref, config_enable_assertion );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_enable_assertion_from_SystemVerilog( config_enable_assertion );
            end
        end
    end

    function automatic void axi_local_set_config_slave_start_addr_from_SystemVerilog( ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param );
        axi_set_config_slave_start_addr_from_SystemVerilog( _interface_ref, config_slave_start_addr );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_slave_start_addr_from_SystemVerilog( config_slave_start_addr );
            end
        end
    end

    function automatic void axi_local_set_config_slave_end_addr_from_SystemVerilog( ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param );
        axi_set_config_slave_end_addr_from_SystemVerilog( _interface_ref, config_slave_end_addr );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_slave_end_addr_from_SystemVerilog( config_slave_end_addr );
            end
        end
    end

    function automatic void axi_local_set_config_support_exclusive_access_from_SystemVerilog( ref bit config_support_exclusive_access_param );
        axi_set_config_support_exclusive_access_from_SystemVerilog( _interface_ref, config_support_exclusive_access );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_support_exclusive_access_from_SystemVerilog( config_support_exclusive_access );
            end
        end
    end

    function automatic void axi_local_set_config_read_data_reordering_depth_from_SystemVerilog( ref int unsigned config_read_data_reordering_depth_param );
        axi_set_config_read_data_reordering_depth_from_SystemVerilog( _interface_ref, config_read_data_reordering_depth );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_read_data_reordering_depth_from_SystemVerilog( config_read_data_reordering_depth );
            end
        end
    end

    function automatic void axi_local_set_config_max_transaction_time_factor_from_SystemVerilog( ref int unsigned config_max_transaction_time_factor_param );
        axi_set_config_max_transaction_time_factor_from_SystemVerilog( _interface_ref, config_max_transaction_time_factor );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_transaction_time_factor_from_SystemVerilog( config_max_transaction_time_factor );
            end
        end
    end

    function automatic void axi_local_set_config_timeout_max_data_transfer_from_SystemVerilog( ref int config_timeout_max_data_transfer_param );
        axi_set_config_timeout_max_data_transfer_from_SystemVerilog( _interface_ref, config_timeout_max_data_transfer );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_timeout_max_data_transfer_from_SystemVerilog( config_timeout_max_data_transfer );
            end
        end
    end

    function automatic void axi_local_set_config_burst_timeout_factor_from_SystemVerilog( ref int unsigned config_burst_timeout_factor_param );
        axi_set_config_burst_timeout_factor_from_SystemVerilog( _interface_ref, config_burst_timeout_factor );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_burst_timeout_factor_from_SystemVerilog( config_burst_timeout_factor );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( ref int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
        axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( _interface_ref, config_max_latency_AWVALID_assertion_to_AWREADY );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( config_max_latency_AWVALID_assertion_to_AWREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( ref int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
        axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( _interface_ref, config_max_latency_ARVALID_assertion_to_ARREADY );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( config_max_latency_ARVALID_assertion_to_ARREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( ref int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
        axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( _interface_ref, config_max_latency_RVALID_assertion_to_RREADY );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( config_max_latency_RVALID_assertion_to_RREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( ref int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
        axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( _interface_ref, config_max_latency_BVALID_assertion_to_BREADY );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( config_max_latency_BVALID_assertion_to_BREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( ref int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
        axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( _interface_ref, config_max_latency_WVALID_assertion_to_WREADY );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( config_max_latency_WVALID_assertion_to_WREADY );
            end
        end
    end

    function automatic void axi_local_set_config_master_error_position_from_SystemVerilog( ref axi_error_e config_master_error_position_param );
        axi_set_config_master_error_position_from_SystemVerilog( _interface_ref, config_master_error_position );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_master_error_position_from_SystemVerilog( config_master_error_position );
            end
        end
    end

    function automatic void axi_local_set_config_setup_time_from_SystemVerilog( ref int config_setup_time_param );
        axi_set_config_setup_time_from_SystemVerilog( _interface_ref, config_setup_time );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_setup_time_from_SystemVerilog( config_setup_time );
            end
        end
    end

    function automatic void axi_local_set_config_hold_time_from_SystemVerilog( ref int config_hold_time_param );
        axi_set_config_hold_time_from_SystemVerilog( _interface_ref, config_hold_time );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_hold_time_from_SystemVerilog( config_hold_time );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_wr_from_SystemVerilog( ref int config_max_outstanding_wr_param );
        axi_set_config_max_outstanding_wr_from_SystemVerilog( _interface_ref, config_max_outstanding_wr );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_wr_from_SystemVerilog( config_max_outstanding_wr );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_rd_from_SystemVerilog( ref int config_max_outstanding_rd_param );
        axi_set_config_max_outstanding_rd_from_SystemVerilog( _interface_ref, config_max_outstanding_rd );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_rd_from_SystemVerilog( config_max_outstanding_rd );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_rw_from_SystemVerilog( ref int config_max_outstanding_rw_param );
        axi_set_config_max_outstanding_rw_from_SystemVerilog( _interface_ref, config_max_outstanding_rw );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_rw_from_SystemVerilog( config_max_outstanding_rw );
            end
        end
    end

    function automatic void axi_local_set_config_is_issuing_from_SystemVerilog( ref bit config_is_issuing_param );
        axi_set_config_is_issuing_from_SystemVerilog( _interface_ref, config_is_issuing );
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_is_issuing_from_SystemVerilog( config_is_issuing );
            end
        end
    end

    //-------------------------------------------------------------------------
    // Transaction interface
    //-------------------------------------------------------------------------

    task automatic dvc_activate_rw_transaction
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp[],
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref axi_rw_e read_or_write,
        ref int address_to_data_latency,
        ref int data_to_response_latency,
        ref int write_address_to_data_delay,
        ref int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        ref int address_valid_delay,
        ref int data_valid_delay[],
        ref int write_response_valid_delay,
        ref int address_ready_delay,
        ref int data_ready_delay[],
        ref int write_response_ready_delay,
        ref bit write_data_with_address,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_valid_delay_DIMS0;
                automatic int data_ready_delay_DIMS0;
            // Call function to provide sized and unsized params.
            // In addition gets back updated sizes of unsized params.
            axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, data_words_DIMS0, write_strobes, write_strobes_DIMS0, resp, resp_DIMS0, addr_user, data_user, data_user_DIMS0, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay, write_data_beats_delay_DIMS0, address_valid_delay, data_valid_delay, data_valid_delay_DIMS0, write_response_valid_delay, address_ready_delay, data_ready_delay, data_ready_delay_DIMS0, write_response_ready_delay, write_data_with_address, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_strobes_DIMS0 != 0)
            begin
                write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                write_strobes = new [1];  // Create dummy instead of a zero sized array
            end
            if (resp_DIMS0 != 0)
            begin
                resp = new [resp_DIMS0];
            end
            else
            begin
                resp = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                write_data_beats_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_valid_delay_DIMS0 != 0)
            begin
                data_valid_delay = new [data_valid_delay_DIMS0];
            end
            else
            begin
                data_valid_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_ready_delay_DIMS0 != 0)
            begin
                data_ready_delay = new [data_ready_delay_DIMS0];
            end
            else
            begin
                data_ready_delay = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, write_strobes, resp, addr_user, data_user, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay, address_valid_delay, data_valid_delay, write_response_valid_delay, address_ready_delay, data_ready_delay, write_response_ready_delay, write_data_with_address, _unit_id); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (write_strobes_DIMS0 == 0)
                write_strobes.delete;  // Delete each zero sized param
            if (resp_DIMS0 == 0)
                resp.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (write_data_beats_delay_DIMS0 == 0)
                write_data_beats_delay.delete;  // Delete each zero sized param
            if (data_valid_delay_DIMS0 == 0)
                data_valid_delay.delete;  // Delete each zero sized param
            if (data_ready_delay_DIMS0 == 0)
                data_ready_delay.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_rw_transaction
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp[],
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output axi_rw_e read_or_write,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        output int address_valid_delay,
        ref int data_valid_delay[],
        output int write_response_valid_delay,
        output int address_ready_delay,
        ref int data_ready_delay[],
        output int write_response_ready_delay,
        output bit write_data_with_address,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_valid_delay_DIMS0;
                automatic int data_ready_delay_DIMS0;
            // Call function to get unsized params sizes.
            axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, resp_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_valid_delay_DIMS0, data_ready_delay_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_strobes_DIMS0 != 0)
            begin
                write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                write_strobes = new [1];  // Create dummy instead of a zero sized array
            end
            if (resp_DIMS0 != 0)
            begin
                resp = new [resp_DIMS0];
            end
            else
            begin
                resp = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                write_data_beats_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_valid_delay_DIMS0 != 0)
            begin
                data_valid_delay = new [data_valid_delay_DIMS0];
            end
            else
            begin
                data_valid_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_ready_delay_DIMS0 != 0)
            begin
                data_ready_delay = new [data_ready_delay_DIMS0];
            end
            else
            begin
                data_ready_delay = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, write_strobes, resp, addr_user, data_user, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay, address_valid_delay, data_valid_delay, write_response_valid_delay, address_ready_delay, data_ready_delay, write_response_ready_delay, write_data_with_address, _unit_id, _using); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (write_strobes_DIMS0 == 0)
                write_strobes.delete;  // Delete each zero sized param
            if (resp_DIMS0 == 0)
                resp.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (write_data_beats_delay_DIMS0 == 0)
                write_data_beats_delay.delete;  // Delete each zero sized param
            if (data_valid_delay_DIMS0 == 0)
                data_valid_delay.delete;  // Delete each zero sized param
            if (data_ready_delay_DIMS0 == 0)
                data_ready_delay.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_AXI_read
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref int address_to_data_latency,
        ref longint addr_start_time,
        ref longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        ref int address_valid_delay,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to provide sized and unsized params.
            // In addition gets back updated sizes of unsized params.
            axi_AXI_read_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, data_words_DIMS0, resp, resp_DIMS0, addr_user, data_user, data_user_DIMS0, address_to_data_latency, addr_start_time, addr_end_time, data_start_time, data_start_time_DIMS0, data_end_time, data_end_time_DIMS0, address_valid_delay, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (resp_DIMS0 != 0)
            begin
                resp = new [resp_DIMS0];
            end
            else
            begin
                resp = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_start_time_DIMS0 != 0)
            begin
                data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                data_start_time = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_end_time_DIMS0 != 0)
            begin
                data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                data_end_time = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, resp, addr_user, data_user, address_to_data_latency, addr_start_time, addr_end_time, data_start_time, data_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (resp_DIMS0 == 0)
                resp.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (data_start_time_DIMS0 == 0)
                data_start_time.delete;  // Delete each zero sized param
            if (data_end_time_DIMS0 == 0)
                data_end_time.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_AXI_read
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output int address_to_data_latency,
        output longint addr_start_time,
        output longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        output int address_valid_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_AXI_read_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, resp_DIMS0, data_user_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (resp_DIMS0 != 0)
            begin
                resp = new [resp_DIMS0];
            end
            else
            begin
                resp = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_start_time_DIMS0 != 0)
            begin
                data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                data_start_time = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_end_time_DIMS0 != 0)
            begin
                data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                data_end_time = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, resp, addr_user, data_user, address_to_data_latency, addr_start_time, addr_end_time, data_start_time, data_end_time, address_valid_delay, _unit_id, _using); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (resp_DIMS0 == 0)
                resp.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (data_start_time_DIMS0 == 0)
                data_start_time.delete;  // Delete each zero sized param
            if (data_end_time_DIMS0 == 0)
                data_end_time.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_AXI_write
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp,
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref int address_to_data_latency,
        ref int data_to_response_latency,
        ref int write_address_to_data_delay,
        ref int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        ref longint addr_start_time,
        ref longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        ref longint wr_resp_start_time,
        ref longint wr_resp_end_time,
        ref int address_valid_delay,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to provide sized and unsized params.
            // In addition gets back updated sizes of unsized params.
            axi_AXI_write_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, data_words_DIMS0, write_strobes, write_strobes_DIMS0, resp, addr_user, data_user, data_user_DIMS0, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay, write_data_beats_delay_DIMS0, addr_start_time, addr_end_time, data_start_time, data_start_time_DIMS0, data_end_time, data_end_time_DIMS0, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_strobes_DIMS0 != 0)
            begin
                write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                write_strobes = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                write_data_beats_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_start_time_DIMS0 != 0)
            begin
                data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                data_start_time = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_end_time_DIMS0 != 0)
            begin
                data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                data_end_time = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, write_strobes, resp, addr_user, data_user, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay, addr_start_time, addr_end_time, data_start_time, data_end_time, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (write_strobes_DIMS0 == 0)
                write_strobes.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (write_data_beats_delay_DIMS0 == 0)
                write_data_beats_delay.delete;  // Delete each zero sized param
            if (data_start_time_DIMS0 == 0)
                data_start_time.delete;  // Delete each zero sized param
            if (data_end_time_DIMS0 == 0)
                data_end_time.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_AXI_write
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output axi_response_e resp,
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        output longint addr_start_time,
        output longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        output longint wr_resp_start_time,
        output longint wr_resp_end_time,
        output int address_valid_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_AXI_write_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_strobes_DIMS0 != 0)
            begin
                write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                write_strobes = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                write_data_beats_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_start_time_DIMS0 != 0)
            begin
                data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                data_start_time = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_end_time_DIMS0 != 0)
            begin
                data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                data_end_time = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, addr, size, burst, lock, cache, prot, id, burst_length, data_words, write_strobes, resp, addr_user, data_user, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay, addr_start_time, addr_end_time, data_start_time, data_end_time, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id, _using); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (write_strobes_DIMS0 == 0)
                write_strobes.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (write_data_beats_delay_DIMS0 == 0)
                write_data_beats_delay.delete;  // Delete each zero sized param
            if (data_start_time_DIMS0 == 0)
                data_start_time.delete;  // Delete each zero sized param
            if (data_end_time_DIMS0 == 0)
                data_end_time.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_data_resp
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref axi_response_e resp,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref longint data_start,
        ref longint data_end,
        ref longint response_start,
        ref int write_data_beats_delay[],
        ref longint data_beat_start_time[],
        ref longint data_beat_end_time[],
        ref longint response_end_time,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_beat_start_time_DIMS0;
                automatic int data_beat_end_time_DIMS0;
            // Call function to provide sized and unsized params.
            // In addition gets back updated sizes of unsized params.
            axi_data_resp_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, data_words, data_words_DIMS0, write_strobes, write_strobes_DIMS0, id, resp, data_user, data_user_DIMS0, resp_user, data_start, data_end, response_start, write_data_beats_delay, write_data_beats_delay_DIMS0, data_beat_start_time, data_beat_start_time_DIMS0, data_beat_end_time, data_beat_end_time_DIMS0, response_end_time, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_strobes_DIMS0 != 0)
            begin
                write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                write_strobes = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                write_data_beats_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_beat_start_time_DIMS0 != 0)
            begin
                data_beat_start_time = new [data_beat_start_time_DIMS0];
            end
            else
            begin
                data_beat_start_time = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_beat_end_time_DIMS0 != 0)
            begin
                data_beat_end_time = new [data_beat_end_time_DIMS0];
            end
            else
            begin
                data_beat_end_time = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, data_words, write_strobes, id, resp, data_user, resp_user, data_start, data_end, response_start, write_data_beats_delay, data_beat_start_time, data_beat_end_time, response_end_time, _unit_id); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (write_strobes_DIMS0 == 0)
                write_strobes.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (write_data_beats_delay_DIMS0 == 0)
                write_data_beats_delay.delete;  // Delete each zero sized param
            if (data_beat_start_time_DIMS0 == 0)
                data_beat_start_time.delete;  // Delete each zero sized param
            if (data_beat_end_time_DIMS0 == 0)
                data_beat_end_time.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_data_resp
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_response_e resp,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output longint data_start,
        output longint data_end,
        output longint response_start,
        ref int write_data_beats_delay[],
        ref longint data_beat_start_time[],
        ref longint data_beat_end_time[],
        output longint response_end_time,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_beat_start_time_DIMS0;
                automatic int data_beat_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_data_resp_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_beat_start_time_DIMS0, data_beat_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_strobes_DIMS0 != 0)
            begin
                write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                write_strobes = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                write_data_beats_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_beat_start_time_DIMS0 != 0)
            begin
                data_beat_start_time = new [data_beat_start_time_DIMS0];
            end
            else
            begin
                data_beat_start_time = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_beat_end_time_DIMS0 != 0)
            begin
                data_beat_end_time = new [data_beat_end_time_DIMS0];
            end
            else
            begin
                data_beat_end_time = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, data_words, write_strobes, id, resp, data_user, resp_user, data_start, data_end, response_start, write_data_beats_delay, data_beat_start_time, data_beat_end_time, response_end_time, _unit_id, _using); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (write_strobes_DIMS0 == 0)
                write_strobes.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (write_data_beats_delay_DIMS0 == 0)
                write_data_beats_delay.delete;  // Delete each zero sized param
            if (data_beat_start_time_DIMS0 == 0)
                data_beat_start_time.delete;  // Delete each zero sized param
            if (data_beat_end_time_DIMS0 == 0)
                data_beat_end_time.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to provide sized and unsized params.
            axi_read_data_burst_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, data_words, resp, id, data_user, data_start_time, data_end_time, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, resp_DIMS0, data_user_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (resp_DIMS0 != 0)
            begin
                resp = new [resp_DIMS0];
            end
            else
            begin
                resp = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_start_time_DIMS0 != 0)
            begin
                data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                data_start_time = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_end_time_DIMS0 != 0)
            begin
                data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                data_end_time = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, data_words, resp, id, data_user, data_start_time, data_end_time, _unit_id, _using); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (resp_DIMS0 == 0)
                resp.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (data_start_time_DIMS0 == 0)
                data_start_time.delete;  // Delete each zero sized param
            if (data_end_time_DIMS0 == 0)
                data_end_time.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref int write_data_beats_delay[],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to provide sized and unsized params.
            axi_write_data_burst_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, data_words, write_strobes, id, data_user, write_data_beats_delay, data_start_time, data_end_time, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref int write_data_beats_delay[],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                data_words = new [data_words_DIMS0];
            end
            else
            begin
                data_words = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_strobes_DIMS0 != 0)
            begin
                write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                write_strobes = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_user_DIMS0 != 0)
            begin
                data_user = new [data_user_DIMS0];
            end
            else
            begin
                data_user = new [1];  // Create dummy instead of a zero sized array
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                write_data_beats_delay = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_start_time_DIMS0 != 0)
            begin
                data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                data_start_time = new [1];  // Create dummy instead of a zero sized array
            end
            if (data_end_time_DIMS0 != 0)
            begin
                data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                data_end_time = new [1];  // Create dummy instead of a zero sized array
            end
            // Call function to get the sized and unsized params
            axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, data_words, write_strobes, id, data_user, write_data_beats_delay, data_start_time, data_end_time, _unit_id, _using); // DPI call to imported task
            if (data_words_DIMS0 == 0)
                data_words.delete;  // Delete each zero sized param
            if (write_strobes_DIMS0 == 0)
                write_strobes.delete;  // Delete each zero sized param
            if (data_user_DIMS0 == 0)
                data_user.delete;  // Delete each zero sized param
            if (write_data_beats_delay_DIMS0 == 0)
                write_data_beats_delay.delete;  // Delete each zero sized param
            if (data_start_time_DIMS0 == 0)
                data_start_time.delete;  // Delete each zero sized param
            if (data_end_time_DIMS0 == 0)
                data_end_time.delete;  // Delete each zero sized param
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, addr, burst_length, size, burst, lock, cache, prot, id, addr_user, address_valid_delay, address_ready_delay, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, addr, burst_length, size, burst, lock, cache, prot, id, addr_user, address_valid_delay, address_ready_delay, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_read_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, data, resp, id, data_user, data_ready_delay, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, last, data, resp, id, data_user, data_ready_delay, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, addr, burst_length, size, burst, lock, cache, prot, id, addr_user, address_valid_delay, address_ready_delay, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, addr, burst_length, size, burst, lock, cache, prot, id, addr_user, address_valid_delay, address_ready_delay, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, data, write_strobes, id, data_user, data_ready_delay, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, last, data, write_strobes, id, data_user, data_ready_delay, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_resp_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int write_response_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, resp, id, resp_user, write_response_ready_delay, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_resp_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        output int write_response_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, resp, id, resp_user, write_response_ready_delay, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_read_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, addr, burst_length, size, burst, lock, cache, prot, id, addr_user, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, addr, burst_length, size, burst, lock, cache, prot, id, addr_user, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_read_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_read_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, data, resp, id, data_user, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, last, data, resp, id, data_user, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_read_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, addr, burst_length, size, burst, lock, cache, prot, id, addr_user, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, addr, burst_length, size, burst, lock, cache, prot, id, addr_user, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, data, strb, id, data_user, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, last, data, strb, id, data_user, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_resp_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, resp, id, resp_user, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_resp_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, resp, id, resp_user, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_resp_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_resp_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask


    //-------------------------------------------------------------------------
    // Generic Interface Configuration Support
    //

    import "DPI-C" context axi_set_interface = function void axi_set_interface
    (
        input int what,
        input int arg1,
        input int arg2,
        input int arg3,
        input int arg4,
        input int arg5,
        input int arg6,
        input int arg7,
        input int arg8,
        input int arg9,
        input int arg10
    );
    import "DPI-C" context axi_get_interface = function int axi_get_interface
    (
        input int what,
        input int arg1,
        input int arg2,
        input int arg3,
        input int arg4,
        input int arg5,
        input int arg6,
        input int arg7,
        input int arg8,
        input int arg9
    );


    //-------------------------------------------------------------------------
    // Functions to get the hierarchic name of this interface
    //
    import "DPI-C" context axi_get_full_name = function string axi_get_full_name();


    //-------------------------------------------------------------------------
    // Abstraction level Support
    //

    import "DPI-C" context axi_set_master_end_abstraction_level =
    function void axi_set_master_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_master_end_abstraction_level =
    function void axi_get_master_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_slave_end_abstraction_level =
    function void axi_set_slave_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_slave_end_abstraction_level =
    function void axi_get_slave_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_clock_source_end_abstraction_level =
    function void axi_set_clock_source_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_clock_source_end_abstraction_level =
    function void axi_get_clock_source_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_reset_source_end_abstraction_level =
    function void axi_set_reset_source_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_reset_source_end_abstraction_level =
    function void axi_get_reset_source_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );

    //-------------------------------------------------------------------------
    // Wire Level Interface Support
    //
    logic internal_ACLK = 'z;
    logic internal_ARESETn = 'z;
    logic internal_AWVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  internal_AWADDR = 'z;
    logic [3:0] internal_AWLEN = 'z;
    logic [2:0] internal_AWSIZE = 'z;
    logic [1:0] internal_AWBURST = 'z;
    logic [1:0] internal_AWLOCK = 'z;
    logic [3:0] internal_AWCACHE = 'z;
    logic [2:0] internal_AWPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_AWID = 'z;
    logic internal_AWREADY = 'z;
    logic [7:0] internal_AWUSER = 'z;
    logic internal_ARVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  internal_ARADDR = 'z;
    logic [3:0] internal_ARLEN = 'z;
    logic [2:0] internal_ARSIZE = 'z;
    logic [1:0] internal_ARBURST = 'z;
    logic [1:0] internal_ARLOCK = 'z;
    logic [3:0] internal_ARCACHE = 'z;
    logic [2:0] internal_ARPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_ARID = 'z;
    logic internal_ARREADY = 'z;
    logic [7:0] internal_ARUSER = 'z;
    logic internal_RVALID = 'z;
    logic internal_RLAST = 'z;
    logic [((AXI_RDATA_WIDTH) - 1):0]  internal_RDATA = 'z;
    logic [1:0] internal_RRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_RID = 'z;
    logic internal_RREADY = 'z;
    logic [7:0] internal_RUSER = 'z;
    logic internal_WVALID = 'z;
    logic internal_WLAST = 'z;
    logic [((AXI_WDATA_WIDTH) - 1):0]  internal_WDATA = 'z;
    logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  internal_WSTRB = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_WID = 'z;
    logic internal_WREADY = 'z;
    logic [7:0] internal_WUSER = 'z;
    logic internal_BVALID = 'z;
    logic [1:0] internal_BRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_BID = 'z;
    logic internal_BREADY = 'z;
    logic [7:0] internal_BUSER = 'z;

    import "DPI-C" context function void axi_set_ACLK_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit ACLK_param
    );
    import "DPI-C" context function void axi_get_ACLK_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit ACLK_param

    );
    export "DPI-C" function axi_initialise_ACLK_from_CY;

    import "DPI-C" context function void axi_set_ARESETn_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARESETn_param
    );
    import "DPI-C" context function void axi_get_ARESETn_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARESETn_param

    );
    export "DPI-C" function axi_initialise_ARESETn_from_CY;

    import "DPI-C" context function void axi_set_AWVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic AWVALID_param
    );
    import "DPI-C" context function void axi_get_AWVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic AWVALID_param

    );
    export "DPI-C" function axi_initialise_AWVALID_from_CY;

    import "DPI-C" context function void axi_set_AWADDR_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_ADDRESS_WIDTH) - 1):0]  AWADDR_param
    );
    import "DPI-C" context function void axi_get_AWADDR_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_ADDRESS_WIDTH) - 1):0]  AWADDR_param

    );
    export "DPI-C" function axi_initialise_AWADDR_from_CY;

    import "DPI-C" context function void axi_set_AWLEN_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] AWLEN_param
    );
    import "DPI-C" context function void axi_get_AWLEN_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] AWLEN_param

    );
    export "DPI-C" function axi_initialise_AWLEN_from_CY;

    import "DPI-C" context function void axi_set_AWSIZE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] AWSIZE_param
    );
    import "DPI-C" context function void axi_get_AWSIZE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] AWSIZE_param

    );
    export "DPI-C" function axi_initialise_AWSIZE_from_CY;

    import "DPI-C" context function void axi_set_AWBURST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] AWBURST_param
    );
    import "DPI-C" context function void axi_get_AWBURST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] AWBURST_param

    );
    export "DPI-C" function axi_initialise_AWBURST_from_CY;

    import "DPI-C" context function void axi_set_AWLOCK_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] AWLOCK_param
    );
    import "DPI-C" context function void axi_get_AWLOCK_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] AWLOCK_param

    );
    export "DPI-C" function axi_initialise_AWLOCK_from_CY;

    import "DPI-C" context function void axi_set_AWCACHE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] AWCACHE_param
    );
    import "DPI-C" context function void axi_get_AWCACHE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] AWCACHE_param

    );
    export "DPI-C" function axi_initialise_AWCACHE_from_CY;

    import "DPI-C" context function void axi_set_AWPROT_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] AWPROT_param
    );
    import "DPI-C" context function void axi_get_AWPROT_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] AWPROT_param

    );
    export "DPI-C" function axi_initialise_AWPROT_from_CY;

    import "DPI-C" context function void axi_set_AWID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_ID_WIDTH) - 1):0]  AWID_param
    );
    import "DPI-C" context function void axi_get_AWID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_ID_WIDTH) - 1):0]  AWID_param

    );
    export "DPI-C" function axi_initialise_AWID_from_CY;

    import "DPI-C" context function void axi_set_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic AWREADY_param
    );
    import "DPI-C" context function void axi_get_AWREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic AWREADY_param

    );
    export "DPI-C" function axi_initialise_AWREADY_from_CY;

    import "DPI-C" context function void axi_set_AWUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] AWUSER_param
    );
    import "DPI-C" context function void axi_get_AWUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] AWUSER_param

    );
    export "DPI-C" function axi_initialise_AWUSER_from_CY;

    import "DPI-C" context function void axi_set_ARVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARVALID_param
    );
    import "DPI-C" context function void axi_get_ARVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARVALID_param

    );
    export "DPI-C" function axi_initialise_ARVALID_from_CY;

    import "DPI-C" context function void axi_set_ARADDR_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_ADDRESS_WIDTH) - 1):0]  ARADDR_param
    );
    import "DPI-C" context function void axi_get_ARADDR_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_ADDRESS_WIDTH) - 1):0]  ARADDR_param

    );
    export "DPI-C" function axi_initialise_ARADDR_from_CY;

    import "DPI-C" context function void axi_set_ARLEN_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] ARLEN_param
    );
    import "DPI-C" context function void axi_get_ARLEN_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] ARLEN_param

    );
    export "DPI-C" function axi_initialise_ARLEN_from_CY;

    import "DPI-C" context function void axi_set_ARSIZE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] ARSIZE_param
    );
    import "DPI-C" context function void axi_get_ARSIZE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] ARSIZE_param

    );
    export "DPI-C" function axi_initialise_ARSIZE_from_CY;

    import "DPI-C" context function void axi_set_ARBURST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] ARBURST_param
    );
    import "DPI-C" context function void axi_get_ARBURST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] ARBURST_param

    );
    export "DPI-C" function axi_initialise_ARBURST_from_CY;

    import "DPI-C" context function void axi_set_ARLOCK_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] ARLOCK_param
    );
    import "DPI-C" context function void axi_get_ARLOCK_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] ARLOCK_param

    );
    export "DPI-C" function axi_initialise_ARLOCK_from_CY;

    import "DPI-C" context function void axi_set_ARCACHE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] ARCACHE_param
    );
    import "DPI-C" context function void axi_get_ARCACHE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] ARCACHE_param

    );
    export "DPI-C" function axi_initialise_ARCACHE_from_CY;

    import "DPI-C" context function void axi_set_ARPROT_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] ARPROT_param
    );
    import "DPI-C" context function void axi_get_ARPROT_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] ARPROT_param

    );
    export "DPI-C" function axi_initialise_ARPROT_from_CY;

    import "DPI-C" context function void axi_set_ARID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_ID_WIDTH) - 1):0]  ARID_param
    );
    import "DPI-C" context function void axi_get_ARID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_ID_WIDTH) - 1):0]  ARID_param

    );
    export "DPI-C" function axi_initialise_ARID_from_CY;

    import "DPI-C" context function void axi_set_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARREADY_param
    );
    import "DPI-C" context function void axi_get_ARREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARREADY_param

    );
    export "DPI-C" function axi_initialise_ARREADY_from_CY;

    import "DPI-C" context function void axi_set_ARUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] ARUSER_param
    );
    import "DPI-C" context function void axi_get_ARUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] ARUSER_param

    );
    export "DPI-C" function axi_initialise_ARUSER_from_CY;

    import "DPI-C" context function void axi_set_RVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RVALID_param
    );
    import "DPI-C" context function void axi_get_RVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RVALID_param

    );
    export "DPI-C" function axi_initialise_RVALID_from_CY;

    import "DPI-C" context function void axi_set_RLAST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RLAST_param
    );
    import "DPI-C" context function void axi_get_RLAST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RLAST_param

    );
    export "DPI-C" function axi_initialise_RLAST_from_CY;

    import "DPI-C" context function void axi_set_RDATA_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_RDATA_WIDTH) - 1):0]  RDATA_param
    );
    import "DPI-C" context function void axi_get_RDATA_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_RDATA_WIDTH) - 1):0]  RDATA_param

    );
    export "DPI-C" function axi_initialise_RDATA_from_CY;

    import "DPI-C" context function void axi_set_RRESP_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] RRESP_param
    );
    import "DPI-C" context function void axi_get_RRESP_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] RRESP_param

    );
    export "DPI-C" function axi_initialise_RRESP_from_CY;

    import "DPI-C" context function void axi_set_RID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_ID_WIDTH) - 1):0]  RID_param
    );
    import "DPI-C" context function void axi_get_RID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_ID_WIDTH) - 1):0]  RID_param

    );
    export "DPI-C" function axi_initialise_RID_from_CY;

    import "DPI-C" context function void axi_set_RREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RREADY_param
    );
    import "DPI-C" context function void axi_get_RREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RREADY_param

    );
    export "DPI-C" function axi_initialise_RREADY_from_CY;

    import "DPI-C" context function void axi_set_RUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] RUSER_param
    );
    import "DPI-C" context function void axi_get_RUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] RUSER_param

    );
    export "DPI-C" function axi_initialise_RUSER_from_CY;

    import "DPI-C" context function void axi_set_WVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WVALID_param
    );
    import "DPI-C" context function void axi_get_WVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WVALID_param

    );
    export "DPI-C" function axi_initialise_WVALID_from_CY;

    import "DPI-C" context function void axi_set_WLAST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WLAST_param
    );
    import "DPI-C" context function void axi_get_WLAST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WLAST_param

    );
    export "DPI-C" function axi_initialise_WLAST_from_CY;

    import "DPI-C" context function void axi_set_WDATA_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_WDATA_WIDTH) - 1):0]  WDATA_param
    );
    import "DPI-C" context function void axi_get_WDATA_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_WDATA_WIDTH) - 1):0]  WDATA_param

    );
    export "DPI-C" function axi_initialise_WDATA_from_CY;

    import "DPI-C" context function void axi_set_WSTRB_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  WSTRB_param
    );
    import "DPI-C" context function void axi_get_WSTRB_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  WSTRB_param

    );
    export "DPI-C" function axi_initialise_WSTRB_from_CY;

    import "DPI-C" context function void axi_set_WID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_ID_WIDTH) - 1):0]  WID_param
    );
    import "DPI-C" context function void axi_get_WID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_ID_WIDTH) - 1):0]  WID_param

    );
    export "DPI-C" function axi_initialise_WID_from_CY;

    import "DPI-C" context function void axi_set_WREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WREADY_param
    );
    import "DPI-C" context function void axi_get_WREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WREADY_param

    );
    export "DPI-C" function axi_initialise_WREADY_from_CY;

    import "DPI-C" context function void axi_set_WUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] WUSER_param
    );
    import "DPI-C" context function void axi_get_WUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] WUSER_param

    );
    export "DPI-C" function axi_initialise_WUSER_from_CY;

    import "DPI-C" context function void axi_set_BVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic BVALID_param
    );
    import "DPI-C" context function void axi_get_BVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic BVALID_param

    );
    export "DPI-C" function axi_initialise_BVALID_from_CY;

    import "DPI-C" context function void axi_set_BRESP_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] BRESP_param
    );
    import "DPI-C" context function void axi_get_BRESP_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] BRESP_param

    );
    export "DPI-C" function axi_initialise_BRESP_from_CY;

    import "DPI-C" context function void axi_set_BID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [((AXI_ID_WIDTH) - 1):0]  BID_param
    );
    import "DPI-C" context function void axi_get_BID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [((AXI_ID_WIDTH) - 1):0]  BID_param

    );
    export "DPI-C" function axi_initialise_BID_from_CY;

    import "DPI-C" context function void axi_set_BREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic BREADY_param
    );
    import "DPI-C" context function void axi_get_BREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic BREADY_param

    );
    export "DPI-C" function axi_initialise_BREADY_from_CY;

    import "DPI-C" context function void axi_set_BUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] BUSER_param
    );
    import "DPI-C" context function void axi_get_BUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] BUSER_param

    );
    export "DPI-C" function axi_initialise_BUSER_from_CY;

    import "DPI-C" context function void axi_set_config_write_ctrl_to_data_mintime_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_write_ctrl_to_data_mintime_param
    );
    import "DPI-C" context function void axi_get_config_write_ctrl_to_data_mintime_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_write_ctrl_to_data_mintime_param

    );
    export "DPI-C" function axi_set_config_write_ctrl_to_data_mintime_from_CY;

    import "DPI-C" context function void axi_set_config_master_write_delay_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_master_write_delay_param
    );
    import "DPI-C" context function void axi_get_deprecated_config_master_write_delay_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_master_write_delay_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_master_write_delay_param

    );
    export "DPI-C" function axi_set_config_master_write_delay_from_CY;

    import "DPI-C" context function void axi_set_config_enable_all_assertions_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_enable_all_assertions_param
    );
    import "DPI-C" context function void axi_get_config_enable_all_assertions_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_enable_all_assertions_param

    );
    export "DPI-C" function axi_set_config_enable_all_assertions_from_CY;

    import "DPI-C" context function void axi_set_config_enable_assertion_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param
    );
    import "DPI-C" context function void axi_get_config_enable_assertion_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param

    );
    export "DPI-C" function axi_set_config_enable_assertion_from_CY;

    import "DPI-C" context function void axi_set_config_slave_start_addr_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param
    );
    import "DPI-C" context function void axi_get_deprecated_config_slave_start_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_slave_start_addr_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param

    );
    export "DPI-C" function axi_set_config_slave_start_addr_from_CY;

    import "DPI-C" context function void axi_set_config_slave_end_addr_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param
    );
    import "DPI-C" context function void axi_get_deprecated_config_slave_end_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_slave_end_addr_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param

    );
    export "DPI-C" function axi_set_config_slave_end_addr_from_CY;

    import "DPI-C" context function void axi_set_config_support_exclusive_access_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_support_exclusive_access_param
    );
    import "DPI-C" context function void axi_get_config_support_exclusive_access_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_support_exclusive_access_param

    );
    export "DPI-C" function axi_set_config_support_exclusive_access_from_CY;

    import "DPI-C" context function void axi_set_config_read_data_reordering_depth_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_read_data_reordering_depth_param
    );
    import "DPI-C" context function void axi_get_config_read_data_reordering_depth_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_read_data_reordering_depth_param

    );
    export "DPI-C" function axi_set_config_read_data_reordering_depth_from_CY;

    import "DPI-C" context function void axi_set_config_max_transaction_time_factor_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_transaction_time_factor_param
    );
    import "DPI-C" context function void axi_get_config_max_transaction_time_factor_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_transaction_time_factor_param

    );
    export "DPI-C" function axi_set_config_max_transaction_time_factor_from_CY;

    import "DPI-C" context function void axi_set_config_timeout_max_data_transfer_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_timeout_max_data_transfer_param
    );
    import "DPI-C" context function void axi_get_config_timeout_max_data_transfer_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_timeout_max_data_transfer_param

    );
    export "DPI-C" function axi_set_config_timeout_max_data_transfer_from_CY;

    import "DPI-C" context function void axi_set_config_burst_timeout_factor_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_burst_timeout_factor_param
    );
    import "DPI-C" context function void axi_get_config_burst_timeout_factor_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_burst_timeout_factor_param

    );
    export "DPI-C" function axi_set_config_burst_timeout_factor_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param
    );
    import "DPI-C" context function void axi_get_config_max_latency_AWVALID_assertion_to_AWREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param
    );
    import "DPI-C" context function void axi_get_config_max_latency_ARVALID_assertion_to_ARREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_RVALID_assertion_to_RREADY_param
    );
    import "DPI-C" context function void axi_get_config_max_latency_RVALID_assertion_to_RREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_RVALID_assertion_to_RREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_BVALID_assertion_to_BREADY_param
    );
    import "DPI-C" context function void axi_get_config_max_latency_BVALID_assertion_to_BREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_BVALID_assertion_to_BREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_WVALID_assertion_to_WREADY_param
    );
    import "DPI-C" context function void axi_get_config_max_latency_WVALID_assertion_to_WREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_WVALID_assertion_to_WREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_CY;

    import "DPI-C" context function void axi_set_config_master_error_position_from_SystemVerilog
    (
        input longint _iface_ref,
        input axi_error_e config_master_error_position_param
    );
    import "DPI-C" context function void axi_get_deprecated_config_master_error_position_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_master_error_position_into_SystemVerilog
    (
        input longint _iface_ref,
        output axi_error_e config_master_error_position_param

    );
    export "DPI-C" function axi_set_config_master_error_position_from_CY;

    import "DPI-C" context function void axi_set_config_setup_time_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_setup_time_param
    );
    import "DPI-C" context function void axi_get_config_setup_time_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_setup_time_param

    );
    export "DPI-C" function axi_set_config_setup_time_from_CY;

    import "DPI-C" context function void axi_set_config_hold_time_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_hold_time_param
    );
    import "DPI-C" context function void axi_get_config_hold_time_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_hold_time_param

    );
    export "DPI-C" function axi_set_config_hold_time_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_wr_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_wr_param
    );
    import "DPI-C" context function void axi_get_config_max_outstanding_wr_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_wr_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_wr_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_rd_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_rd_param
    );
    import "DPI-C" context function void axi_get_config_max_outstanding_rd_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_rd_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_rd_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_rw_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_rw_param
    );
    import "DPI-C" context function void axi_get_config_max_outstanding_rw_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_rw_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_rw_from_CY;

    import "DPI-C" context function void axi_set_config_is_issuing_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_is_issuing_param
    );
    import "DPI-C" context function void axi_get_config_is_issuing_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_is_issuing_param

    );
    export "DPI-C" function axi_set_config_is_issuing_from_CY;

    function void axi_initialise_ACLK_from_CY();
        internal_ACLK = 'z;
        m_ACLK = 'z;
    endfunction

    function void axi_initialise_ARESETn_from_CY();
        internal_ARESETn = 'z;
        m_ARESETn = 'z;
    endfunction

    function void axi_initialise_AWVALID_from_CY();
        internal_AWVALID = 'z;
        m_AWVALID = 'z;
    endfunction

    function void axi_initialise_AWADDR_from_CY();
        internal_AWADDR = 'z;
        m_AWADDR = 'z;
    endfunction

    function void axi_initialise_AWLEN_from_CY();
        internal_AWLEN = 'z;
        m_AWLEN = 'z;
    endfunction

    function void axi_initialise_AWSIZE_from_CY();
        internal_AWSIZE = 'z;
        m_AWSIZE = 'z;
    endfunction

    function void axi_initialise_AWBURST_from_CY();
        internal_AWBURST = 'z;
        m_AWBURST = 'z;
    endfunction

    function void axi_initialise_AWLOCK_from_CY();
        internal_AWLOCK = 'z;
        m_AWLOCK = 'z;
    endfunction

    function void axi_initialise_AWCACHE_from_CY();
        internal_AWCACHE = 'z;
        m_AWCACHE = 'z;
    endfunction

    function void axi_initialise_AWPROT_from_CY();
        internal_AWPROT = 'z;
        m_AWPROT = 'z;
    endfunction

    function void axi_initialise_AWID_from_CY();
        internal_AWID = 'z;
        m_AWID = 'z;
    endfunction

    function void axi_initialise_AWREADY_from_CY();
        internal_AWREADY = 'z;
        m_AWREADY = 'z;
    endfunction

    function void axi_initialise_AWUSER_from_CY();
        internal_AWUSER = 'z;
        m_AWUSER = 'z;
    endfunction

    function void axi_initialise_ARVALID_from_CY();
        internal_ARVALID = 'z;
        m_ARVALID = 'z;
    endfunction

    function void axi_initialise_ARADDR_from_CY();
        internal_ARADDR = 'z;
        m_ARADDR = 'z;
    endfunction

    function void axi_initialise_ARLEN_from_CY();
        internal_ARLEN = 'z;
        m_ARLEN = 'z;
    endfunction

    function void axi_initialise_ARSIZE_from_CY();
        internal_ARSIZE = 'z;
        m_ARSIZE = 'z;
    endfunction

    function void axi_initialise_ARBURST_from_CY();
        internal_ARBURST = 'z;
        m_ARBURST = 'z;
    endfunction

    function void axi_initialise_ARLOCK_from_CY();
        internal_ARLOCK = 'z;
        m_ARLOCK = 'z;
    endfunction

    function void axi_initialise_ARCACHE_from_CY();
        internal_ARCACHE = 'z;
        m_ARCACHE = 'z;
    endfunction

    function void axi_initialise_ARPROT_from_CY();
        internal_ARPROT = 'z;
        m_ARPROT = 'z;
    endfunction

    function void axi_initialise_ARID_from_CY();
        internal_ARID = 'z;
        m_ARID = 'z;
    endfunction

    function void axi_initialise_ARREADY_from_CY();
        internal_ARREADY = 'z;
        m_ARREADY = 'z;
    endfunction

    function void axi_initialise_ARUSER_from_CY();
        internal_ARUSER = 'z;
        m_ARUSER = 'z;
    endfunction

    function void axi_initialise_RVALID_from_CY();
        internal_RVALID = 'z;
        m_RVALID = 'z;
    endfunction

    function void axi_initialise_RLAST_from_CY();
        internal_RLAST = 'z;
        m_RLAST = 'z;
    endfunction

    function void axi_initialise_RDATA_from_CY();
        internal_RDATA = 'z;
        m_RDATA = 'z;
    endfunction

    function void axi_initialise_RRESP_from_CY();
        internal_RRESP = 'z;
        m_RRESP = 'z;
    endfunction

    function void axi_initialise_RID_from_CY();
        internal_RID = 'z;
        m_RID = 'z;
    endfunction

    function void axi_initialise_RREADY_from_CY();
        internal_RREADY = 'z;
        m_RREADY = 'z;
    endfunction

    function void axi_initialise_RUSER_from_CY();
        internal_RUSER = 'z;
        m_RUSER = 'z;
    endfunction

    function void axi_initialise_WVALID_from_CY();
        internal_WVALID = 'z;
        m_WVALID = 'z;
    endfunction

    function void axi_initialise_WLAST_from_CY();
        internal_WLAST = 'z;
        m_WLAST = 'z;
    endfunction

    function void axi_initialise_WDATA_from_CY();
        internal_WDATA = 'z;
        m_WDATA = 'z;
    endfunction

    function void axi_initialise_WSTRB_from_CY();
        internal_WSTRB = 'z;
        m_WSTRB = 'z;
    endfunction

    function void axi_initialise_WID_from_CY();
        internal_WID = 'z;
        m_WID = 'z;
    endfunction

    function void axi_initialise_WREADY_from_CY();
        internal_WREADY = 'z;
        m_WREADY = 'z;
    endfunction

    function void axi_initialise_WUSER_from_CY();
        internal_WUSER = 'z;
        m_WUSER = 'z;
    endfunction

    function void axi_initialise_BVALID_from_CY();
        internal_BVALID = 'z;
        m_BVALID = 'z;
    endfunction

    function void axi_initialise_BRESP_from_CY();
        internal_BRESP = 'z;
        m_BRESP = 'z;
    endfunction

    function void axi_initialise_BID_from_CY();
        internal_BID = 'z;
        m_BID = 'z;
    endfunction

    function void axi_initialise_BREADY_from_CY();
        internal_BREADY = 'z;
        m_BREADY = 'z;
    endfunction

    function void axi_initialise_BUSER_from_CY();
        internal_BUSER = 'z;
        m_BUSER = 'z;
    endfunction

    function void axi_set_config_write_ctrl_to_data_mintime_from_CY( int unsigned config_write_ctrl_to_data_mintime_param );
        config_write_ctrl_to_data_mintime = config_write_ctrl_to_data_mintime_param;
    endfunction

    function void axi_set_config_master_write_delay_from_CY( bit config_master_write_delay_param );
        config_master_write_delay = config_master_write_delay_param;
    endfunction

    function void axi_set_config_enable_all_assertions_from_CY( bit config_enable_all_assertions_param );
        config_enable_all_assertions = config_enable_all_assertions_param;
    endfunction

    function void axi_set_config_enable_assertion_from_CY( bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
        config_enable_assertion = config_enable_assertion_param;
    endfunction

    function void axi_set_config_slave_start_addr_from_CY( bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param );
        config_slave_start_addr = config_slave_start_addr_param;
    endfunction

    function void axi_set_config_slave_end_addr_from_CY( bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param );
        config_slave_end_addr = config_slave_end_addr_param;
    endfunction

    function void axi_set_config_support_exclusive_access_from_CY( bit config_support_exclusive_access_param );
        config_support_exclusive_access = config_support_exclusive_access_param;
    endfunction

    function void axi_set_config_read_data_reordering_depth_from_CY( int unsigned config_read_data_reordering_depth_param );
        config_read_data_reordering_depth = config_read_data_reordering_depth_param;
    endfunction

    function void axi_set_config_max_transaction_time_factor_from_CY( int unsigned config_max_transaction_time_factor_param );
        config_max_transaction_time_factor = config_max_transaction_time_factor_param;
    endfunction

    function void axi_set_config_timeout_max_data_transfer_from_CY( int config_timeout_max_data_transfer_param );
        config_timeout_max_data_transfer = config_timeout_max_data_transfer_param;
    endfunction

    function void axi_set_config_burst_timeout_factor_from_CY( int unsigned config_burst_timeout_factor_param );
        config_burst_timeout_factor = config_burst_timeout_factor_param;
    endfunction

    function void axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_CY( int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
        config_max_latency_AWVALID_assertion_to_AWREADY = config_max_latency_AWVALID_assertion_to_AWREADY_param;
    endfunction

    function void axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_CY( int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
        config_max_latency_ARVALID_assertion_to_ARREADY = config_max_latency_ARVALID_assertion_to_ARREADY_param;
    endfunction

    function void axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_CY( int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
        config_max_latency_RVALID_assertion_to_RREADY = config_max_latency_RVALID_assertion_to_RREADY_param;
    endfunction

    function void axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_CY( int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
        config_max_latency_BVALID_assertion_to_BREADY = config_max_latency_BVALID_assertion_to_BREADY_param;
    endfunction

    function void axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_CY( int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
        config_max_latency_WVALID_assertion_to_WREADY = config_max_latency_WVALID_assertion_to_WREADY_param;
    endfunction

    function void axi_set_config_master_error_position_from_CY( axi_error_e config_master_error_position_param );
        config_master_error_position = config_master_error_position_param;
    endfunction

    function void axi_set_config_setup_time_from_CY( int config_setup_time_param );
        config_setup_time = config_setup_time_param;
    endfunction

    function void axi_set_config_hold_time_from_CY( int config_hold_time_param );
        config_hold_time = config_hold_time_param;
    endfunction

    function void axi_set_config_max_outstanding_wr_from_CY( int config_max_outstanding_wr_param );
        config_max_outstanding_wr = config_max_outstanding_wr_param;
    endfunction

    function void axi_set_config_max_outstanding_rd_from_CY( int config_max_outstanding_rd_param );
        config_max_outstanding_rd = config_max_outstanding_rd_param;
    endfunction

    function void axi_set_config_max_outstanding_rw_from_CY( int config_max_outstanding_rw_param );
        config_max_outstanding_rw = config_max_outstanding_rw_param;
    endfunction

    function void axi_set_config_is_issuing_from_CY( bit config_is_issuing_param );
        config_is_issuing = config_is_issuing_param;
    endfunction



    //--------------------------------------------------------------------------
    //
    // Group:- TLM Interface Support
    //
    //--------------------------------------------------------------------------
    import "DPI-C" context axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog =
    task axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        input bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        input axi_response_e resp[],
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] addr_user,
        input bit [7:0] data_user [],
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout axi_rw_e read_or_write,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        input int write_data_beats_delay[],
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_valid_delay,
        input int data_valid_delay[],
        inout int data_valid_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_response_valid_delay,
        inout int address_ready_delay,
        input int data_ready_delay[],
        inout int data_ready_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_response_ready_delay,
        inout bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        inout bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout axi_response_e resp[],
        inout bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout axi_rw_e read_or_write,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int write_data_beats_delay[],
        inout int address_valid_delay,
        inout int data_valid_delay[],
        inout int write_response_valid_delay,
        inout int address_ready_delay,
        inout int data_ready_delay[],
        inout int write_response_ready_delay,
        inout bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_START_ActivatesActivatingActivate_SystemVerilog =
    function int axi_rw_transaction_START_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        input bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        input axi_response_e resp[],
        inout bit [7:0] addr_user,
        input bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout axi_rw_e read_or_write,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        input int write_data_beats_delay[],
        inout int address_valid_delay,
        input int data_valid_delay[],
        inout int write_response_valid_delay,
        inout int address_ready_delay,
        input int data_ready_delay[],
        inout int write_response_ready_delay,
        inout bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_END_ActivatesActivatingActivate_SystemVerilog =
    function int axi_rw_transaction_END_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_valid_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_ready_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_END_ActivatesActivatingActivate_open_SystemVerilog =
    function int axi_rw_transaction_END_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        inout bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout axi_response_e resp[],
        inout bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout axi_rw_e read_or_write,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int write_data_beats_delay[],
        inout int address_valid_delay,
        inout int data_valid_delay[],
        inout int write_response_valid_delay,
        inout int address_ready_delay,
        inout int data_ready_delay[],
        inout int write_response_ready_delay,
        inout bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog =
    task axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_valid_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_ready_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        inout bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout axi_response_e resp[],
        output bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output axi_rw_e read_or_write,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        inout int write_data_beats_delay[],
        output int address_valid_delay,
        inout int data_valid_delay[],
        output int write_response_valid_delay,
        output int address_ready_delay,
        inout int data_ready_delay[],
        output int write_response_ready_delay,
        output bit write_data_with_address,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_rw_transaction_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_rw_transaction_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_rw_transaction_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_rw_transaction_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_valid_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_ready_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_END_ReceivedReceivingReceive_open_SystemVerilog =
    function int axi_rw_transaction_END_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        inout bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout axi_response_e resp[],
        output bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output axi_rw_e read_or_write,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        inout int write_data_beats_delay[],
        output int address_valid_delay,
        inout int data_valid_delay[],
        output int write_response_valid_delay,
        output int address_ready_delay,
        inout int data_ready_delay[],
        output int write_response_ready_delay,
        output bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_ActivatesActivatingActivate_SystemVerilog =
    task axi_AXI_read_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        input bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        input axi_response_e resp[],
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] addr_user,
        input bit [7:0] data_user [],
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_to_data_latency,
        inout longint addr_start_time,
        inout longint addr_end_time,
        input longint data_start_time[],
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input longint data_end_time[],
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        inout bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        inout axi_response_e resp[],
        inout bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        inout int address_to_data_latency,
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout longint data_start_time[],
        inout longint data_end_time[],
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_START_ActivatesActivatingActivate_SystemVerilog =
    function int axi_AXI_read_START_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        input bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        input axi_response_e resp[],
        inout bit [7:0] addr_user,
        input bit [7:0] data_user [],
        inout int address_to_data_latency,
        inout longint addr_start_time,
        inout longint addr_end_time,
        input longint data_start_time[],
        input longint data_end_time[],
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_END_ActivatesActivatingActivate_SystemVerilog =
    function int axi_AXI_read_END_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_END_ActivatesActivatingActivate_open_SystemVerilog =
    function int axi_AXI_read_END_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        inout bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        inout axi_response_e resp[],
        inout bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        inout int address_to_data_latency,
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout longint data_start_time[],
        inout longint data_end_time[],
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_ReceivedReceivingReceive_SystemVerilog =
    task axi_AXI_read_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        inout bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        inout axi_response_e resp[],
        output bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        output int address_to_data_latency,
        output longint addr_start_time,
        output longint addr_end_time,
        inout longint data_start_time[],
        inout longint data_end_time[],
        output int address_valid_delay,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_read_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_AXI_read_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_read_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_AXI_read_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_END_ReceivedReceivingReceive_open_SystemVerilog =
    function int axi_AXI_read_END_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        inout bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        inout axi_response_e resp[],
        output bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        output int address_to_data_latency,
        output longint addr_start_time,
        output longint addr_end_time,
        inout longint data_start_time[],
        inout longint data_end_time[],
        output int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_ActivatesActivatingActivate_SystemVerilog =
    task axi_AXI_write_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        input bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout axi_response_e resp,
        inout bit [7:0] addr_user,
        input bit [7:0] data_user [],
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        input int write_data_beats_delay[],
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint addr_start_time,
        inout longint addr_end_time,
        input longint data_start_time[],
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input longint data_end_time[],
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint wr_resp_start_time,
        inout longint wr_resp_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout axi_response_e resp,
        inout bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int write_data_beats_delay[],
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout longint data_start_time[],
        inout longint data_end_time[],
        inout longint wr_resp_start_time,
        inout longint wr_resp_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_START_ActivatesActivatingActivate_SystemVerilog =
    function int axi_AXI_write_START_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        input bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout axi_response_e resp,
        inout bit [7:0] addr_user,
        input bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        input int write_data_beats_delay[],
        inout longint addr_start_time,
        inout longint addr_end_time,
        input longint data_start_time[],
        input longint data_end_time[],
        inout longint wr_resp_start_time,
        inout longint wr_resp_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_END_ActivatesActivatingActivate_SystemVerilog =
    function int axi_AXI_write_END_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_END_ActivatesActivatingActivate_open_SystemVerilog =
    function int axi_AXI_write_END_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [3:0] burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout axi_response_e resp,
        inout bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int write_data_beats_delay[],
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout longint data_start_time[],
        inout longint data_end_time[],
        inout longint wr_resp_start_time,
        inout longint wr_resp_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_ReceivedReceivingReceive_SystemVerilog =
    task axi_AXI_write_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output axi_response_e resp,
        output bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        inout int write_data_beats_delay[],
        output longint addr_start_time,
        output longint addr_end_time,
        inout longint data_start_time[],
        inout longint data_end_time[],
        output longint wr_resp_start_time,
        output longint wr_resp_end_time,
        output int address_valid_delay,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_write_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_AXI_write_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_write_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_AXI_write_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_END_ReceivedReceivingReceive_open_SystemVerilog =
    function int axi_AXI_write_END_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output axi_response_e resp,
        output bit [7:0] addr_user,
        inout bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        inout int write_data_beats_delay[],
        output longint addr_start_time,
        output longint addr_end_time,
        inout longint data_start_time[],
        inout longint data_end_time[],
        output longint wr_resp_start_time,
        output longint wr_resp_end_time,
        output int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_ActivatesActivatingActivate_SystemVerilog =
    task axi_data_resp_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int burst_length,
        input bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout axi_response_e resp,
        input bit [7:0] data_user [],
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout longint data_start,
        inout longint data_end,
        inout longint response_start,
        input int write_data_beats_delay[],
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        input longint data_beat_start_time[],
        inout int data_beat_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input longint data_beat_end_time[],
        inout int data_beat_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout axi_response_e resp,
        inout bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout longint data_start,
        inout longint data_end,
        inout longint response_start,
        inout int write_data_beats_delay[],
        inout longint data_beat_start_time[],
        inout longint data_beat_end_time[],
        inout longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_START_ActivatesActivatingActivate_SystemVerilog =
    function int axi_data_resp_START_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        inout int burst_length,
        input bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout axi_response_e resp,
        input bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout longint data_start,
        inout longint data_end,
        inout longint response_start,
        input int write_data_beats_delay[],
        input longint data_beat_start_time[],
        input longint data_beat_end_time[],
        inout longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_END_ActivatesActivatingActivate_SystemVerilog =
    function int axi_data_resp_END_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_END_ActivatesActivatingActivate_open_SystemVerilog =
    function int axi_data_resp_END_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        inout bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout axi_response_e resp,
        inout bit [7:0] data_user [],
        inout bit [7:0] resp_user,
        inout longint data_start,
        inout longint data_end,
        inout longint response_start,
        inout int write_data_beats_delay[],
        inout longint data_beat_start_time[],
        inout longint data_beat_end_time[],
        inout longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_ReceivedReceivingReceive_SystemVerilog =
    task axi_data_resp_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output int burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_response_e resp,
        inout bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output longint data_start,
        output longint data_end,
        output longint response_start,
        inout int write_data_beats_delay[],
        inout longint data_beat_start_time[],
        inout longint data_beat_end_time[],
        output longint response_end_time,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_data_resp_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_data_resp_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_data_resp_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_data_resp_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_END_ReceivedReceivingReceive_open_SystemVerilog =
    function int axi_data_resp_END_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output int burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_response_e resp,
        inout bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output longint data_start,
        output longint data_end,
        output longint response_start,
        inout int write_data_beats_delay[],
        inout longint data_beat_start_time[],
        inout longint data_beat_end_time[],
        output longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_read_data_burst_SendSendingSent_SystemVerilog =
    task axi_read_data_burst_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        input axi_response_e resp[],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user [],
        input longint data_start_time[],
        input longint data_end_time[],
        input int _unit_id
    );
    import "DPI-C" context axi_read_data_burst_START_SendSendingSent_SystemVerilog =
    function int axi_read_data_burst_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        input axi_response_e resp[],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user [],
        input longint data_start_time[],
        input longint data_end_time[],
        input int _unit_id
    );
    import "DPI-C" context axi_read_data_burst_END_SendSendingSent_SystemVerilog =
    function int axi_read_data_burst_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [3:0] burst_length,
        inout bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        inout axi_response_e resp[],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [7:0] data_user [],
        inout longint data_start_time[],
        inout longint data_end_time[],
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_data_burst_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_data_burst_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_data_burst_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_data_burst_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_read_data_burst_END_ReceivedReceivingReceive_open_SystemVerilog =
    function int axi_read_data_burst_END_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [3:0] burst_length,
        inout bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        inout axi_response_e resp[],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [7:0] data_user [],
        inout longint data_start_time[],
        inout longint data_end_time[],
        input int _unit_id
    );
    import "DPI-C" context axi_write_data_burst_SendSendingSent_SystemVerilog =
    task axi_write_data_burst_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int burst_length,
        input bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user [],
        input int write_data_beats_delay[],
        input longint data_start_time[],
        input longint data_end_time[],
        input int _unit_id
    );
    import "DPI-C" context axi_write_data_burst_START_SendSendingSent_SystemVerilog =
    function int axi_write_data_burst_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int burst_length,
        input bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user [],
        input int write_data_beats_delay[],
        input longint data_start_time[],
        input longint data_end_time[],
        input int _unit_id
    );
    import "DPI-C" context axi_write_data_burst_END_SendSendingSent_SystemVerilog =
    function int axi_write_data_burst_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output int burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [7:0] data_user [],
        inout int write_data_beats_delay[],
        inout longint data_start_time[],
        inout longint data_end_time[],
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_data_burst_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_data_burst_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_data_burst_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_data_burst_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_write_data_burst_END_ReceivedReceivingReceive_open_SystemVerilog =
    function int axi_write_data_burst_END_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output int burst_length,
        inout bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        inout bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        inout bit [7:0] data_user [],
        inout int write_data_beats_delay[],
        inout longint data_start_time[],
        inout longint data_end_time[],
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_phase_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_phase_START_SendSendingSent_SystemVerilog =
    function int axi_read_addr_channel_phase_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_phase_END_SendSendingSent_SystemVerilog =
    function int axi_read_addr_channel_phase_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_phase_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_addr_channel_phase_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_phase_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_addr_channel_phase_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_phase_SendSendingSent_SystemVerilog =
    task axi_read_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_phase_START_SendSendingSent_SystemVerilog =
    function int axi_read_channel_phase_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_phase_END_SendSendingSent_SystemVerilog =
    function int axi_read_channel_phase_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_phase_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_channel_phase_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_phase_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_channel_phase_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_phase_START_SendSendingSent_SystemVerilog =
    function int axi_write_addr_channel_phase_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_phase_END_SendSendingSent_SystemVerilog =
    function int axi_write_addr_channel_phase_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_phase_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_addr_channel_phase_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_phase_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_addr_channel_phase_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_phase_START_SendSendingSent_SystemVerilog =
    function int axi_write_channel_phase_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_phase_END_SendSendingSent_SystemVerilog =
    function int axi_write_channel_phase_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_phase_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_channel_phase_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_phase_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_channel_phase_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int write_response_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_phase_START_SendSendingSent_SystemVerilog =
    function int axi_write_resp_channel_phase_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int write_response_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_phase_END_SendSendingSent_SystemVerilog =
    function int axi_write_resp_channel_phase_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        output int write_response_ready_delay,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_phase_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_resp_channel_phase_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_phase_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_resp_channel_phase_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        output int write_response_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_cycle_START_SendSendingSent_SystemVerilog =
    function int axi_read_addr_channel_cycle_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_cycle_END_SendSendingSent_SystemVerilog =
    function int axi_read_addr_channel_cycle_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_addr_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_addr_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_ready_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_ready_START_SendSendingSent_SystemVerilog =
    function int axi_read_addr_channel_ready_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_ready_END_SendSendingSent_SystemVerilog =
    function int axi_read_addr_channel_ready_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_ready_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_addr_channel_ready_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_ready_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_addr_channel_ready_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_read_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_cycle_START_SendSendingSent_SystemVerilog =
    function int axi_read_channel_cycle_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_cycle_END_SendSendingSent_SystemVerilog =
    function int axi_read_channel_cycle_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_ready_SendSendingSent_SystemVerilog =
    task axi_read_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_ready_START_SendSendingSent_SystemVerilog =
    function int axi_read_channel_ready_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_ready_END_SendSendingSent_SystemVerilog =
    function int axi_read_channel_ready_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_ready_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_channel_ready_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_ready_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_read_channel_ready_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_cycle_START_SendSendingSent_SystemVerilog =
    function int axi_write_addr_channel_cycle_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_cycle_END_SendSendingSent_SystemVerilog =
    function int axi_write_addr_channel_cycle_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_addr_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_addr_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_ready_START_SendSendingSent_SystemVerilog =
    function int axi_write_addr_channel_ready_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_ready_END_SendSendingSent_SystemVerilog =
    function int axi_write_addr_channel_ready_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_ready_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_addr_channel_ready_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_ready_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_addr_channel_ready_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_cycle_START_SendSendingSent_SystemVerilog =
    function int axi_write_channel_cycle_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_cycle_END_SendSendingSent_SystemVerilog =
    function int axi_write_channel_cycle_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_ready_START_SendSendingSent_SystemVerilog =
    function int axi_write_channel_ready_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_ready_END_SendSendingSent_SystemVerilog =
    function int axi_write_channel_ready_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_ready_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_channel_ready_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_ready_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_channel_ready_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_cycle_START_SendSendingSent_SystemVerilog =
    function int axi_write_resp_channel_cycle_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_cycle_END_SendSendingSent_SystemVerilog =
    function int axi_write_resp_channel_cycle_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_resp_channel_cycle_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_resp_channel_cycle_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_ready_START_SendSendingSent_SystemVerilog =
    function int axi_write_resp_channel_ready_START_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_ready_END_SendSendingSent_SystemVerilog =
    function int axi_write_resp_channel_ready_END_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_ready_START_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_resp_channel_ready_START_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_ready_END_ReceivedReceivingReceive_SystemVerilog =
    function int axi_write_resp_channel_ready_END_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_fn_rd_txn_valid_lanes = function void fn_rd_txn_valid_lanes_C
    (
        inout bit [((AXI_RDATA_WIDTH / 8) - 1):0] valid_lanes []
    );

    import "DPI-C" context axi_fn_get_wdata_phase_info = function void fn_get_wdata_phase_info_C
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit wdata_last,
        inout bit waddr_rcvd,
        output bit [3:0] burst_length,
        output int beat_num,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  beat_addr
    );

    import "DPI-C" context axi_fn_get_wresp_phase_info = function void fn_get_wresp_phase_info_C
    (
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  wresp_corr_addr
    );

    import "DPI-C" context axi_fn_get_rdata_phase_info = function void fn_get_rdata_phase_info_C
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit rdata_last,
        output bit [3:0] burst_length,
        output int beat_num,
        output bit [((AXI_RDATA_WIDTH / 8) - 1):0]  beat_strobes,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  beat_addr,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  txn_addr
    );

    import "DPI-C" context axi_fn_get_max_os_per_id = function void fn_get_max_os_per_id_C
    (
        output int max_waddr_os,
        output int max_wdata_os
    );

    import "DPI-C" context axi_get_rw_txns_in_prog = function void get_rw_txns_in_prog_C
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_rw_txn_counts_s txn_counts
    );

    import "DPI-C" context axi_fn_add_addr_map_entry = function void fn_add_addr_map_entry_C
    (
        input string region,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input longint unsigned size
    );

    import "DPI-C" context axi_fn_add_wr_delay = function void fn_add_wr_delay_C
    (
        input string region,
        input bit [17:0] id,
        input int unsigned addr2data,
        input int unsigned data2data[]
    );

    import "DPI-C" context axi_fn_delete_wr_delay = function void fn_delete_wr_delay_C
    (
        input string region,
        input bit [17:0] id
    );

    import "DPI-C" context axi_fn_set_wr_def_delays = function void fn_set_wr_def_delays_C
    (
        input int unsigned min_addr2data,
        input int unsigned min_data2data[],
        input int unsigned max_addr2data,
        input int unsigned max_data2data[]
    );

    // Waiter task and control
    reg wait_for_control = 0;

    always @(posedge wait_for_control)
    begin
        disable wait_for;
        wait_for_control = 0;
    end

    export "DPI-C" axi_wait_for = task wait_for;

    task wait_for();
        begin
            wait(0 == 1);
        end
    endtask

    // Drive wires (from Cohesive) 
    assign ACLK = internal_ACLK;
    assign ARESETn = internal_ARESETn;
    assign AWVALID = internal_AWVALID;
    assign AWADDR = internal_AWADDR;
    assign AWLEN = internal_AWLEN;
    assign AWSIZE = internal_AWSIZE;
    assign AWBURST = internal_AWBURST;
    assign AWLOCK = internal_AWLOCK;
    assign AWCACHE = internal_AWCACHE;
    assign AWPROT = internal_AWPROT;
    assign AWID = internal_AWID;
    assign AWREADY = internal_AWREADY;
    assign AWUSER = internal_AWUSER;
    assign ARVALID = internal_ARVALID;
    assign ARADDR = internal_ARADDR;
    assign ARLEN = internal_ARLEN;
    assign ARSIZE = internal_ARSIZE;
    assign ARBURST = internal_ARBURST;
    assign ARLOCK = internal_ARLOCK;
    assign ARCACHE = internal_ARCACHE;
    assign ARPROT = internal_ARPROT;
    assign ARID = internal_ARID;
    assign ARREADY = internal_ARREADY;
    assign ARUSER = internal_ARUSER;
    assign RVALID = internal_RVALID;
    assign RLAST = internal_RLAST;
    assign RDATA = internal_RDATA;
    assign RRESP = internal_RRESP;
    assign RID = internal_RID;
    assign RREADY = internal_RREADY;
    assign RUSER = internal_RUSER;
    assign WVALID = internal_WVALID;
    assign WLAST = internal_WLAST;
    assign WDATA = internal_WDATA;
    assign WSTRB = internal_WSTRB;
    assign WID = internal_WID;
    assign WREADY = internal_WREADY;
    assign WUSER = internal_WUSER;
    assign BVALID = internal_BVALID;
    assign BRESP = internal_BRESP;
    assign BID = internal_BID;
    assign BREADY = internal_BREADY;
    assign BUSER = internal_BUSER;
    // Drive wires (from User) 
    assign ACLK = m_ACLK;
    assign ARESETn = m_ARESETn;
    assign AWVALID = m_AWVALID;
    assign AWADDR = m_AWADDR;
    assign AWLEN = m_AWLEN;
    assign AWSIZE = m_AWSIZE;
    assign AWBURST = m_AWBURST;
    assign AWLOCK = m_AWLOCK;
    assign AWCACHE = m_AWCACHE;
    assign AWPROT = m_AWPROT;
    assign AWID = m_AWID;
    assign AWREADY = m_AWREADY;
    assign AWUSER = m_AWUSER;
    assign ARVALID = m_ARVALID;
    assign ARADDR = m_ARADDR;
    assign ARLEN = m_ARLEN;
    assign ARSIZE = m_ARSIZE;
    assign ARBURST = m_ARBURST;
    assign ARLOCK = m_ARLOCK;
    assign ARCACHE = m_ARCACHE;
    assign ARPROT = m_ARPROT;
    assign ARID = m_ARID;
    assign ARREADY = m_ARREADY;
    assign ARUSER = m_ARUSER;
    assign RVALID = m_RVALID;
    assign RLAST = m_RLAST;
    assign RDATA = m_RDATA;
    assign RRESP = m_RRESP;
    assign RID = m_RID;
    assign RREADY = m_RREADY;
    assign RUSER = m_RUSER;
    assign WVALID = m_WVALID;
    assign WLAST = m_WLAST;
    assign WDATA = m_WDATA;
    assign WSTRB = m_WSTRB;
    assign WID = m_WID;
    assign WREADY = m_WREADY;
    assign WUSER = m_WUSER;
    assign BVALID = m_BVALID;
    assign BRESP = m_BRESP;
    assign BID = m_BID;
    assign BREADY = m_BREADY;
    assign BUSER = m_BUSER;

    reg ACLK_changed = 0;
    reg ARESETn_changed = 0;
    reg AWVALID_changed = 0;
    reg AWADDR_changed = 0;
    reg AWLEN_changed = 0;
    reg AWSIZE_changed = 0;
    reg AWBURST_changed = 0;
    reg AWLOCK_changed = 0;
    reg AWCACHE_changed = 0;
    reg AWPROT_changed = 0;
    reg AWID_changed = 0;
    reg AWREADY_changed = 0;
    reg AWUSER_changed = 0;
    reg ARVALID_changed = 0;
    reg ARADDR_changed = 0;
    reg ARLEN_changed = 0;
    reg ARSIZE_changed = 0;
    reg ARBURST_changed = 0;
    reg ARLOCK_changed = 0;
    reg ARCACHE_changed = 0;
    reg ARPROT_changed = 0;
    reg ARID_changed = 0;
    reg ARREADY_changed = 0;
    reg ARUSER_changed = 0;
    reg RVALID_changed = 0;
    reg RLAST_changed = 0;
    reg RDATA_changed = 0;
    reg RRESP_changed = 0;
    reg RID_changed = 0;
    reg RREADY_changed = 0;
    reg RUSER_changed = 0;
    reg WVALID_changed = 0;
    reg WLAST_changed = 0;
    reg WDATA_changed = 0;
    reg WSTRB_changed = 0;
    reg WID_changed = 0;
    reg WREADY_changed = 0;
    reg WUSER_changed = 0;
    reg BVALID_changed = 0;
    reg BRESP_changed = 0;
    reg BID_changed = 0;
    reg BREADY_changed = 0;
    reg BUSER_changed = 0;
    reg config_write_ctrl_to_data_mintime_changed = 0;
    reg config_master_write_delay_changed = 0;
    reg config_enable_all_assertions_changed = 0;
    reg config_enable_assertion_changed = 0;
    reg config_slave_start_addr_changed = 0;
    reg config_slave_end_addr_changed = 0;
    reg config_support_exclusive_access_changed = 0;
    reg config_read_data_reordering_depth_changed = 0;
    reg config_max_transaction_time_factor_changed = 0;
    reg config_timeout_max_data_transfer_changed = 0;
    reg config_burst_timeout_factor_changed = 0;
    reg config_max_latency_AWVALID_assertion_to_AWREADY_changed = 0;
    reg config_max_latency_ARVALID_assertion_to_ARREADY_changed = 0;
    reg config_max_latency_RVALID_assertion_to_RREADY_changed = 0;
    reg config_max_latency_BVALID_assertion_to_BREADY_changed = 0;
    reg config_max_latency_WVALID_assertion_to_WREADY_changed = 0;
    reg config_master_error_position_changed = 0;
    reg config_setup_time_changed = 0;
    reg config_hold_time_changed = 0;
    reg config_max_outstanding_wr_changed = 0;
    reg config_max_outstanding_rd_changed = 0;
    reg config_max_outstanding_rw_changed = 0;
    reg config_is_issuing_changed = 0;
    // Timeless transaction monitor
    reg timeless_trans_control= 0;

    // SV wire change monitors

    always @( ACLK or posedge _check_t0_values )
    begin
        axi_set_ACLK_from_SystemVerilog(_interface_ref, ACLK); // DPI call to imported task
    end

    always @( ARESETn or posedge _check_t0_values )
    begin
        axi_set_ARESETn_from_SystemVerilog(_interface_ref, ARESETn); // DPI call to imported task
    end

    always @( AWVALID or posedge _check_t0_values )
    begin
        axi_set_AWVALID_from_SystemVerilog(_interface_ref, AWVALID); // DPI call to imported task
    end

    always @( AWADDR or posedge _check_t0_values )
    begin
        axi_set_AWADDR_from_SystemVerilog(_interface_ref, AWADDR); // DPI call to imported task
    end

    always @( AWLEN or posedge _check_t0_values )
    begin
        axi_set_AWLEN_from_SystemVerilog(_interface_ref, AWLEN); // DPI call to imported task
    end

    always @( AWSIZE or posedge _check_t0_values )
    begin
        axi_set_AWSIZE_from_SystemVerilog(_interface_ref, AWSIZE); // DPI call to imported task
    end

    always @( AWBURST or posedge _check_t0_values )
    begin
        axi_set_AWBURST_from_SystemVerilog(_interface_ref, AWBURST); // DPI call to imported task
    end

    always @( AWLOCK or posedge _check_t0_values )
    begin
        axi_set_AWLOCK_from_SystemVerilog(_interface_ref, AWLOCK); // DPI call to imported task
    end

    always @( AWCACHE or posedge _check_t0_values )
    begin
        axi_set_AWCACHE_from_SystemVerilog(_interface_ref, AWCACHE); // DPI call to imported task
    end

    always @( AWPROT or posedge _check_t0_values )
    begin
        axi_set_AWPROT_from_SystemVerilog(_interface_ref, AWPROT); // DPI call to imported task
    end

    always @( AWID or posedge _check_t0_values )
    begin
        axi_set_AWID_from_SystemVerilog(_interface_ref, AWID); // DPI call to imported task
    end

    always @( AWREADY or posedge _check_t0_values )
    begin
        axi_set_AWREADY_from_SystemVerilog(_interface_ref, AWREADY); // DPI call to imported task
    end

    always @( AWUSER or posedge _check_t0_values )
    begin
        axi_set_AWUSER_from_SystemVerilog(_interface_ref, AWUSER); // DPI call to imported task
    end

    always @( ARVALID or posedge _check_t0_values )
    begin
        axi_set_ARVALID_from_SystemVerilog(_interface_ref, ARVALID); // DPI call to imported task
    end

    always @( ARADDR or posedge _check_t0_values )
    begin
        axi_set_ARADDR_from_SystemVerilog(_interface_ref, ARADDR); // DPI call to imported task
    end

    always @( ARLEN or posedge _check_t0_values )
    begin
        axi_set_ARLEN_from_SystemVerilog(_interface_ref, ARLEN); // DPI call to imported task
    end

    always @( ARSIZE or posedge _check_t0_values )
    begin
        axi_set_ARSIZE_from_SystemVerilog(_interface_ref, ARSIZE); // DPI call to imported task
    end

    always @( ARBURST or posedge _check_t0_values )
    begin
        axi_set_ARBURST_from_SystemVerilog(_interface_ref, ARBURST); // DPI call to imported task
    end

    always @( ARLOCK or posedge _check_t0_values )
    begin
        axi_set_ARLOCK_from_SystemVerilog(_interface_ref, ARLOCK); // DPI call to imported task
    end

    always @( ARCACHE or posedge _check_t0_values )
    begin
        axi_set_ARCACHE_from_SystemVerilog(_interface_ref, ARCACHE); // DPI call to imported task
    end

    always @( ARPROT or posedge _check_t0_values )
    begin
        axi_set_ARPROT_from_SystemVerilog(_interface_ref, ARPROT); // DPI call to imported task
    end

    always @( ARID or posedge _check_t0_values )
    begin
        axi_set_ARID_from_SystemVerilog(_interface_ref, ARID); // DPI call to imported task
    end

    always @( ARREADY or posedge _check_t0_values )
    begin
        axi_set_ARREADY_from_SystemVerilog(_interface_ref, ARREADY); // DPI call to imported task
    end

    always @( ARUSER or posedge _check_t0_values )
    begin
        axi_set_ARUSER_from_SystemVerilog(_interface_ref, ARUSER); // DPI call to imported task
    end

    always @( RVALID or posedge _check_t0_values )
    begin
        axi_set_RVALID_from_SystemVerilog(_interface_ref, RVALID); // DPI call to imported task
    end

    always @( RLAST or posedge _check_t0_values )
    begin
        axi_set_RLAST_from_SystemVerilog(_interface_ref, RLAST); // DPI call to imported task
    end

    always @( RDATA or posedge _check_t0_values )
    begin
        axi_set_RDATA_from_SystemVerilog(_interface_ref, RDATA); // DPI call to imported task
    end

    always @( RRESP or posedge _check_t0_values )
    begin
        axi_set_RRESP_from_SystemVerilog(_interface_ref, RRESP); // DPI call to imported task
    end

    always @( RID or posedge _check_t0_values )
    begin
        axi_set_RID_from_SystemVerilog(_interface_ref, RID); // DPI call to imported task
    end

    always @( RREADY or posedge _check_t0_values )
    begin
        axi_set_RREADY_from_SystemVerilog(_interface_ref, RREADY); // DPI call to imported task
    end

    always @( RUSER or posedge _check_t0_values )
    begin
        axi_set_RUSER_from_SystemVerilog(_interface_ref, RUSER); // DPI call to imported task
    end

    always @( WVALID or posedge _check_t0_values )
    begin
        axi_set_WVALID_from_SystemVerilog(_interface_ref, WVALID); // DPI call to imported task
    end

    always @( WLAST or posedge _check_t0_values )
    begin
        axi_set_WLAST_from_SystemVerilog(_interface_ref, WLAST); // DPI call to imported task
    end

    always @( WDATA or posedge _check_t0_values )
    begin
        axi_set_WDATA_from_SystemVerilog(_interface_ref, WDATA); // DPI call to imported task
    end

    always @( WSTRB or posedge _check_t0_values )
    begin
        axi_set_WSTRB_from_SystemVerilog(_interface_ref, WSTRB); // DPI call to imported task
    end

    always @( WID or posedge _check_t0_values )
    begin
        axi_set_WID_from_SystemVerilog(_interface_ref, WID); // DPI call to imported task
    end

    always @( WREADY or posedge _check_t0_values )
    begin
        axi_set_WREADY_from_SystemVerilog(_interface_ref, WREADY); // DPI call to imported task
    end

    always @( WUSER or posedge _check_t0_values )
    begin
        axi_set_WUSER_from_SystemVerilog(_interface_ref, WUSER); // DPI call to imported task
    end

    always @( BVALID or posedge _check_t0_values )
    begin
        axi_set_BVALID_from_SystemVerilog(_interface_ref, BVALID); // DPI call to imported task
    end

    always @( BRESP or posedge _check_t0_values )
    begin
        axi_set_BRESP_from_SystemVerilog(_interface_ref, BRESP); // DPI call to imported task
    end

    always @( BID or posedge _check_t0_values )
    begin
        axi_set_BID_from_SystemVerilog(_interface_ref, BID); // DPI call to imported task
    end

    always @( BREADY or posedge _check_t0_values )
    begin
        axi_set_BREADY_from_SystemVerilog(_interface_ref, BREADY); // DPI call to imported task
    end

    always @( BUSER or posedge _check_t0_values )
    begin
        axi_set_BUSER_from_SystemVerilog(_interface_ref, BUSER); // DPI call to imported task
    end


    // CY wire and variable changed flag monitors

    always @(posedge ACLK_changed or posedge _check_t0_values )
    begin
        while (ACLK_changed == 1'b1)
        begin
            axi_get_ACLK_into_SystemVerilog( _interface_ref, internal_ACLK ); // DPI call to imported task
            ACLK_changed = 1'b0;
            #0 if ( ACLK !== internal_ACLK )
            begin
                axi_set_ACLK_from_SystemVerilog( _interface_ref, ACLK );
            end
        end
    end

    always @(posedge ARESETn_changed or posedge _check_t0_values )
    begin
        while (ARESETn_changed == 1'b1)
        begin
            axi_get_ARESETn_into_SystemVerilog( _interface_ref, internal_ARESETn ); // DPI call to imported task
            ARESETn_changed = 1'b0;
            #0 if ( ARESETn !== internal_ARESETn )
            begin
                axi_set_ARESETn_from_SystemVerilog( _interface_ref, ARESETn );
            end
        end
    end

    always @(posedge AWVALID_changed or posedge _check_t0_values )
    begin
        while (AWVALID_changed == 1'b1)
        begin
            axi_get_AWVALID_into_SystemVerilog( _interface_ref, internal_AWVALID ); // DPI call to imported task
            AWVALID_changed = 1'b0;
            #0 if ( AWVALID !== internal_AWVALID )
            begin
                axi_set_AWVALID_from_SystemVerilog( _interface_ref, AWVALID );
            end
        end
    end

    always @(posedge AWADDR_changed or posedge _check_t0_values )
    begin
        while (AWADDR_changed == 1'b1)
        begin
            axi_get_AWADDR_into_SystemVerilog( _interface_ref, internal_AWADDR ); // DPI call to imported task
            AWADDR_changed = 1'b0;
            #0 if ( AWADDR !== internal_AWADDR )
            begin
                axi_set_AWADDR_from_SystemVerilog( _interface_ref, AWADDR );
            end
        end
    end

    always @(posedge AWLEN_changed or posedge _check_t0_values )
    begin
        while (AWLEN_changed == 1'b1)
        begin
            axi_get_AWLEN_into_SystemVerilog( _interface_ref, internal_AWLEN ); // DPI call to imported task
            AWLEN_changed = 1'b0;
            #0 if ( AWLEN !== internal_AWLEN )
            begin
                axi_set_AWLEN_from_SystemVerilog( _interface_ref, AWLEN );
            end
        end
    end

    always @(posedge AWSIZE_changed or posedge _check_t0_values )
    begin
        while (AWSIZE_changed == 1'b1)
        begin
            axi_get_AWSIZE_into_SystemVerilog( _interface_ref, internal_AWSIZE ); // DPI call to imported task
            AWSIZE_changed = 1'b0;
            #0 if ( AWSIZE !== internal_AWSIZE )
            begin
                axi_set_AWSIZE_from_SystemVerilog( _interface_ref, AWSIZE );
            end
        end
    end

    always @(posedge AWBURST_changed or posedge _check_t0_values )
    begin
        while (AWBURST_changed == 1'b1)
        begin
            axi_get_AWBURST_into_SystemVerilog( _interface_ref, internal_AWBURST ); // DPI call to imported task
            AWBURST_changed = 1'b0;
            #0 if ( AWBURST !== internal_AWBURST )
            begin
                axi_set_AWBURST_from_SystemVerilog( _interface_ref, AWBURST );
            end
        end
    end

    always @(posedge AWLOCK_changed or posedge _check_t0_values )
    begin
        while (AWLOCK_changed == 1'b1)
        begin
            axi_get_AWLOCK_into_SystemVerilog( _interface_ref, internal_AWLOCK ); // DPI call to imported task
            AWLOCK_changed = 1'b0;
            #0 if ( AWLOCK !== internal_AWLOCK )
            begin
                axi_set_AWLOCK_from_SystemVerilog( _interface_ref, AWLOCK );
            end
        end
    end

    always @(posedge AWCACHE_changed or posedge _check_t0_values )
    begin
        while (AWCACHE_changed == 1'b1)
        begin
            axi_get_AWCACHE_into_SystemVerilog( _interface_ref, internal_AWCACHE ); // DPI call to imported task
            AWCACHE_changed = 1'b0;
            #0 if ( AWCACHE !== internal_AWCACHE )
            begin
                axi_set_AWCACHE_from_SystemVerilog( _interface_ref, AWCACHE );
            end
        end
    end

    always @(posedge AWPROT_changed or posedge _check_t0_values )
    begin
        while (AWPROT_changed == 1'b1)
        begin
            axi_get_AWPROT_into_SystemVerilog( _interface_ref, internal_AWPROT ); // DPI call to imported task
            AWPROT_changed = 1'b0;
            #0 if ( AWPROT !== internal_AWPROT )
            begin
                axi_set_AWPROT_from_SystemVerilog( _interface_ref, AWPROT );
            end
        end
    end

    always @(posedge AWID_changed or posedge _check_t0_values )
    begin
        while (AWID_changed == 1'b1)
        begin
            axi_get_AWID_into_SystemVerilog( _interface_ref, internal_AWID ); // DPI call to imported task
            AWID_changed = 1'b0;
            #0 if ( AWID !== internal_AWID )
            begin
                axi_set_AWID_from_SystemVerilog( _interface_ref, AWID );
            end
        end
    end

    always @(posedge AWREADY_changed or posedge _check_t0_values )
    begin
        while (AWREADY_changed == 1'b1)
        begin
            axi_get_AWREADY_into_SystemVerilog( _interface_ref, internal_AWREADY ); // DPI call to imported task
            AWREADY_changed = 1'b0;
            #0 if ( AWREADY !== internal_AWREADY )
            begin
                axi_set_AWREADY_from_SystemVerilog( _interface_ref, AWREADY );
            end
        end
    end

    always @(posedge AWUSER_changed or posedge _check_t0_values )
    begin
        while (AWUSER_changed == 1'b1)
        begin
            axi_get_AWUSER_into_SystemVerilog( _interface_ref, internal_AWUSER ); // DPI call to imported task
            AWUSER_changed = 1'b0;
            #0 if ( AWUSER !== internal_AWUSER )
            begin
                axi_set_AWUSER_from_SystemVerilog( _interface_ref, AWUSER );
            end
        end
    end

    always @(posedge ARVALID_changed or posedge _check_t0_values )
    begin
        while (ARVALID_changed == 1'b1)
        begin
            axi_get_ARVALID_into_SystemVerilog( _interface_ref, internal_ARVALID ); // DPI call to imported task
            ARVALID_changed = 1'b0;
            #0 if ( ARVALID !== internal_ARVALID )
            begin
                axi_set_ARVALID_from_SystemVerilog( _interface_ref, ARVALID );
            end
        end
    end

    always @(posedge ARADDR_changed or posedge _check_t0_values )
    begin
        while (ARADDR_changed == 1'b1)
        begin
            axi_get_ARADDR_into_SystemVerilog( _interface_ref, internal_ARADDR ); // DPI call to imported task
            ARADDR_changed = 1'b0;
            #0 if ( ARADDR !== internal_ARADDR )
            begin
                axi_set_ARADDR_from_SystemVerilog( _interface_ref, ARADDR );
            end
        end
    end

    always @(posedge ARLEN_changed or posedge _check_t0_values )
    begin
        while (ARLEN_changed == 1'b1)
        begin
            axi_get_ARLEN_into_SystemVerilog( _interface_ref, internal_ARLEN ); // DPI call to imported task
            ARLEN_changed = 1'b0;
            #0 if ( ARLEN !== internal_ARLEN )
            begin
                axi_set_ARLEN_from_SystemVerilog( _interface_ref, ARLEN );
            end
        end
    end

    always @(posedge ARSIZE_changed or posedge _check_t0_values )
    begin
        while (ARSIZE_changed == 1'b1)
        begin
            axi_get_ARSIZE_into_SystemVerilog( _interface_ref, internal_ARSIZE ); // DPI call to imported task
            ARSIZE_changed = 1'b0;
            #0 if ( ARSIZE !== internal_ARSIZE )
            begin
                axi_set_ARSIZE_from_SystemVerilog( _interface_ref, ARSIZE );
            end
        end
    end

    always @(posedge ARBURST_changed or posedge _check_t0_values )
    begin
        while (ARBURST_changed == 1'b1)
        begin
            axi_get_ARBURST_into_SystemVerilog( _interface_ref, internal_ARBURST ); // DPI call to imported task
            ARBURST_changed = 1'b0;
            #0 if ( ARBURST !== internal_ARBURST )
            begin
                axi_set_ARBURST_from_SystemVerilog( _interface_ref, ARBURST );
            end
        end
    end

    always @(posedge ARLOCK_changed or posedge _check_t0_values )
    begin
        while (ARLOCK_changed == 1'b1)
        begin
            axi_get_ARLOCK_into_SystemVerilog( _interface_ref, internal_ARLOCK ); // DPI call to imported task
            ARLOCK_changed = 1'b0;
            #0 if ( ARLOCK !== internal_ARLOCK )
            begin
                axi_set_ARLOCK_from_SystemVerilog( _interface_ref, ARLOCK );
            end
        end
    end

    always @(posedge ARCACHE_changed or posedge _check_t0_values )
    begin
        while (ARCACHE_changed == 1'b1)
        begin
            axi_get_ARCACHE_into_SystemVerilog( _interface_ref, internal_ARCACHE ); // DPI call to imported task
            ARCACHE_changed = 1'b0;
            #0 if ( ARCACHE !== internal_ARCACHE )
            begin
                axi_set_ARCACHE_from_SystemVerilog( _interface_ref, ARCACHE );
            end
        end
    end

    always @(posedge ARPROT_changed or posedge _check_t0_values )
    begin
        while (ARPROT_changed == 1'b1)
        begin
            axi_get_ARPROT_into_SystemVerilog( _interface_ref, internal_ARPROT ); // DPI call to imported task
            ARPROT_changed = 1'b0;
            #0 if ( ARPROT !== internal_ARPROT )
            begin
                axi_set_ARPROT_from_SystemVerilog( _interface_ref, ARPROT );
            end
        end
    end

    always @(posedge ARID_changed or posedge _check_t0_values )
    begin
        while (ARID_changed == 1'b1)
        begin
            axi_get_ARID_into_SystemVerilog( _interface_ref, internal_ARID ); // DPI call to imported task
            ARID_changed = 1'b0;
            #0 if ( ARID !== internal_ARID )
            begin
                axi_set_ARID_from_SystemVerilog( _interface_ref, ARID );
            end
        end
    end

    always @(posedge ARREADY_changed or posedge _check_t0_values )
    begin
        while (ARREADY_changed == 1'b1)
        begin
            axi_get_ARREADY_into_SystemVerilog( _interface_ref, internal_ARREADY ); // DPI call to imported task
            ARREADY_changed = 1'b0;
            #0 if ( ARREADY !== internal_ARREADY )
            begin
                axi_set_ARREADY_from_SystemVerilog( _interface_ref, ARREADY );
            end
        end
    end

    always @(posedge ARUSER_changed or posedge _check_t0_values )
    begin
        while (ARUSER_changed == 1'b1)
        begin
            axi_get_ARUSER_into_SystemVerilog( _interface_ref, internal_ARUSER ); // DPI call to imported task
            ARUSER_changed = 1'b0;
            #0 if ( ARUSER !== internal_ARUSER )
            begin
                axi_set_ARUSER_from_SystemVerilog( _interface_ref, ARUSER );
            end
        end
    end

    always @(posedge RVALID_changed or posedge _check_t0_values )
    begin
        while (RVALID_changed == 1'b1)
        begin
            axi_get_RVALID_into_SystemVerilog( _interface_ref, internal_RVALID ); // DPI call to imported task
            RVALID_changed = 1'b0;
            #0 if ( RVALID !== internal_RVALID )
            begin
                axi_set_RVALID_from_SystemVerilog( _interface_ref, RVALID );
            end
        end
    end

    always @(posedge RLAST_changed or posedge _check_t0_values )
    begin
        while (RLAST_changed == 1'b1)
        begin
            axi_get_RLAST_into_SystemVerilog( _interface_ref, internal_RLAST ); // DPI call to imported task
            RLAST_changed = 1'b0;
            #0 if ( RLAST !== internal_RLAST )
            begin
                axi_set_RLAST_from_SystemVerilog( _interface_ref, RLAST );
            end
        end
    end

    always @(posedge RDATA_changed or posedge _check_t0_values )
    begin
        while (RDATA_changed == 1'b1)
        begin
            axi_get_RDATA_into_SystemVerilog( _interface_ref, internal_RDATA ); // DPI call to imported task
            RDATA_changed = 1'b0;
            #0 if ( RDATA !== internal_RDATA )
            begin
                axi_set_RDATA_from_SystemVerilog( _interface_ref, RDATA );
            end
        end
    end

    always @(posedge RRESP_changed or posedge _check_t0_values )
    begin
        while (RRESP_changed == 1'b1)
        begin
            axi_get_RRESP_into_SystemVerilog( _interface_ref, internal_RRESP ); // DPI call to imported task
            RRESP_changed = 1'b0;
            #0 if ( RRESP !== internal_RRESP )
            begin
                axi_set_RRESP_from_SystemVerilog( _interface_ref, RRESP );
            end
        end
    end

    always @(posedge RID_changed or posedge _check_t0_values )
    begin
        while (RID_changed == 1'b1)
        begin
            axi_get_RID_into_SystemVerilog( _interface_ref, internal_RID ); // DPI call to imported task
            RID_changed = 1'b0;
            #0 if ( RID !== internal_RID )
            begin
                axi_set_RID_from_SystemVerilog( _interface_ref, RID );
            end
        end
    end

    always @(posedge RREADY_changed or posedge _check_t0_values )
    begin
        while (RREADY_changed == 1'b1)
        begin
            axi_get_RREADY_into_SystemVerilog( _interface_ref, internal_RREADY ); // DPI call to imported task
            RREADY_changed = 1'b0;
            #0 if ( RREADY !== internal_RREADY )
            begin
                axi_set_RREADY_from_SystemVerilog( _interface_ref, RREADY );
            end
        end
    end

    always @(posedge RUSER_changed or posedge _check_t0_values )
    begin
        while (RUSER_changed == 1'b1)
        begin
            axi_get_RUSER_into_SystemVerilog( _interface_ref, internal_RUSER ); // DPI call to imported task
            RUSER_changed = 1'b0;
            #0 if ( RUSER !== internal_RUSER )
            begin
                axi_set_RUSER_from_SystemVerilog( _interface_ref, RUSER );
            end
        end
    end

    always @(posedge WVALID_changed or posedge _check_t0_values )
    begin
        while (WVALID_changed == 1'b1)
        begin
            axi_get_WVALID_into_SystemVerilog( _interface_ref, internal_WVALID ); // DPI call to imported task
            WVALID_changed = 1'b0;
            #0 if ( WVALID !== internal_WVALID )
            begin
                axi_set_WVALID_from_SystemVerilog( _interface_ref, WVALID );
            end
        end
    end

    always @(posedge WLAST_changed or posedge _check_t0_values )
    begin
        while (WLAST_changed == 1'b1)
        begin
            axi_get_WLAST_into_SystemVerilog( _interface_ref, internal_WLAST ); // DPI call to imported task
            WLAST_changed = 1'b0;
            #0 if ( WLAST !== internal_WLAST )
            begin
                axi_set_WLAST_from_SystemVerilog( _interface_ref, WLAST );
            end
        end
    end

    always @(posedge WDATA_changed or posedge _check_t0_values )
    begin
        while (WDATA_changed == 1'b1)
        begin
            axi_get_WDATA_into_SystemVerilog( _interface_ref, internal_WDATA ); // DPI call to imported task
            WDATA_changed = 1'b0;
            #0 if ( WDATA !== internal_WDATA )
            begin
                axi_set_WDATA_from_SystemVerilog( _interface_ref, WDATA );
            end
        end
    end

    always @(posedge WSTRB_changed or posedge _check_t0_values )
    begin
        while (WSTRB_changed == 1'b1)
        begin
            axi_get_WSTRB_into_SystemVerilog( _interface_ref, internal_WSTRB ); // DPI call to imported task
            WSTRB_changed = 1'b0;
            #0 if ( WSTRB !== internal_WSTRB )
            begin
                axi_set_WSTRB_from_SystemVerilog( _interface_ref, WSTRB );
            end
        end
    end

    always @(posedge WID_changed or posedge _check_t0_values )
    begin
        while (WID_changed == 1'b1)
        begin
            axi_get_WID_into_SystemVerilog( _interface_ref, internal_WID ); // DPI call to imported task
            WID_changed = 1'b0;
            #0 if ( WID !== internal_WID )
            begin
                axi_set_WID_from_SystemVerilog( _interface_ref, WID );
            end
        end
    end

    always @(posedge WREADY_changed or posedge _check_t0_values )
    begin
        while (WREADY_changed == 1'b1)
        begin
            axi_get_WREADY_into_SystemVerilog( _interface_ref, internal_WREADY ); // DPI call to imported task
            WREADY_changed = 1'b0;
            #0 if ( WREADY !== internal_WREADY )
            begin
                axi_set_WREADY_from_SystemVerilog( _interface_ref, WREADY );
            end
        end
    end

    always @(posedge WUSER_changed or posedge _check_t0_values )
    begin
        while (WUSER_changed == 1'b1)
        begin
            axi_get_WUSER_into_SystemVerilog( _interface_ref, internal_WUSER ); // DPI call to imported task
            WUSER_changed = 1'b0;
            #0 if ( WUSER !== internal_WUSER )
            begin
                axi_set_WUSER_from_SystemVerilog( _interface_ref, WUSER );
            end
        end
    end

    always @(posedge BVALID_changed or posedge _check_t0_values )
    begin
        while (BVALID_changed == 1'b1)
        begin
            axi_get_BVALID_into_SystemVerilog( _interface_ref, internal_BVALID ); // DPI call to imported task
            BVALID_changed = 1'b0;
            #0 if ( BVALID !== internal_BVALID )
            begin
                axi_set_BVALID_from_SystemVerilog( _interface_ref, BVALID );
            end
        end
    end

    always @(posedge BRESP_changed or posedge _check_t0_values )
    begin
        while (BRESP_changed == 1'b1)
        begin
            axi_get_BRESP_into_SystemVerilog( _interface_ref, internal_BRESP ); // DPI call to imported task
            BRESP_changed = 1'b0;
            #0 if ( BRESP !== internal_BRESP )
            begin
                axi_set_BRESP_from_SystemVerilog( _interface_ref, BRESP );
            end
        end
    end

    always @(posedge BID_changed or posedge _check_t0_values )
    begin
        while (BID_changed == 1'b1)
        begin
            axi_get_BID_into_SystemVerilog( _interface_ref, internal_BID ); // DPI call to imported task
            BID_changed = 1'b0;
            #0 if ( BID !== internal_BID )
            begin
                axi_set_BID_from_SystemVerilog( _interface_ref, BID );
            end
        end
    end

    always @(posedge BREADY_changed or posedge _check_t0_values )
    begin
        while (BREADY_changed == 1'b1)
        begin
            axi_get_BREADY_into_SystemVerilog( _interface_ref, internal_BREADY ); // DPI call to imported task
            BREADY_changed = 1'b0;
            #0 if ( BREADY !== internal_BREADY )
            begin
                axi_set_BREADY_from_SystemVerilog( _interface_ref, BREADY );
            end
        end
    end

    always @(posedge BUSER_changed or posedge _check_t0_values )
    begin
        while (BUSER_changed == 1'b1)
        begin
            axi_get_BUSER_into_SystemVerilog( _interface_ref, internal_BUSER ); // DPI call to imported task
            BUSER_changed = 1'b0;
            #0 if ( BUSER !== internal_BUSER )
            begin
                axi_set_BUSER_from_SystemVerilog( _interface_ref, BUSER );
            end
        end
    end

    always @(posedge config_write_ctrl_to_data_mintime_changed or posedge _check_t0_values )
    begin
        if (config_write_ctrl_to_data_mintime_changed == 1'b1)
        begin
            axi_get_config_write_ctrl_to_data_mintime_into_SystemVerilog( _interface_ref, config_write_ctrl_to_data_mintime ); // DPI call to imported task
            config_write_ctrl_to_data_mintime_changed = 1'b0;
        end
    end

    always @(posedge config_master_write_delay_changed or posedge _check_t0_values )
    begin
        if (config_master_write_delay_changed == 1'b1)
        begin
            axi_get_config_master_write_delay_into_SystemVerilog( _interface_ref, config_master_write_delay ); // DPI call to imported task
            config_master_write_delay_changed = 1'b0;
        end
    end

    always @(posedge config_enable_all_assertions_changed or posedge _check_t0_values )
    begin
        if (config_enable_all_assertions_changed == 1'b1)
        begin
            axi_get_config_enable_all_assertions_into_SystemVerilog( _interface_ref, config_enable_all_assertions ); // DPI call to imported task
            config_enable_all_assertions_changed = 1'b0;
        end
    end

    always @(posedge config_enable_assertion_changed or posedge _check_t0_values )
    begin
        if (config_enable_assertion_changed == 1'b1)
        begin
            axi_get_config_enable_assertion_into_SystemVerilog( _interface_ref, config_enable_assertion ); // DPI call to imported task
            config_enable_assertion_changed = 1'b0;
        end
    end

    always @(posedge config_slave_start_addr_changed or posedge _check_t0_values )
    begin
        if (config_slave_start_addr_changed == 1'b1)
        begin
            axi_get_config_slave_start_addr_into_SystemVerilog( _interface_ref, config_slave_start_addr ); // DPI call to imported task
            config_slave_start_addr_changed = 1'b0;
        end
    end

    always @(posedge config_slave_end_addr_changed or posedge _check_t0_values )
    begin
        if (config_slave_end_addr_changed == 1'b1)
        begin
            axi_get_config_slave_end_addr_into_SystemVerilog( _interface_ref, config_slave_end_addr ); // DPI call to imported task
            config_slave_end_addr_changed = 1'b0;
        end
    end

    always @(posedge config_support_exclusive_access_changed or posedge _check_t0_values )
    begin
        if (config_support_exclusive_access_changed == 1'b1)
        begin
            axi_get_config_support_exclusive_access_into_SystemVerilog( _interface_ref, config_support_exclusive_access ); // DPI call to imported task
            config_support_exclusive_access_changed = 1'b0;
        end
    end

    always @(posedge config_read_data_reordering_depth_changed or posedge _check_t0_values )
    begin
        if (config_read_data_reordering_depth_changed == 1'b1)
        begin
            axi_get_config_read_data_reordering_depth_into_SystemVerilog( _interface_ref, config_read_data_reordering_depth ); // DPI call to imported task
            config_read_data_reordering_depth_changed = 1'b0;
        end
    end

    always @(posedge config_max_transaction_time_factor_changed or posedge _check_t0_values )
    begin
        if (config_max_transaction_time_factor_changed == 1'b1)
        begin
            axi_get_config_max_transaction_time_factor_into_SystemVerilog( _interface_ref, config_max_transaction_time_factor ); // DPI call to imported task
            config_max_transaction_time_factor_changed = 1'b0;
        end
    end

    always @(posedge config_timeout_max_data_transfer_changed or posedge _check_t0_values )
    begin
        if (config_timeout_max_data_transfer_changed == 1'b1)
        begin
            axi_get_config_timeout_max_data_transfer_into_SystemVerilog( _interface_ref, config_timeout_max_data_transfer ); // DPI call to imported task
            config_timeout_max_data_transfer_changed = 1'b0;
        end
    end

    always @(posedge config_burst_timeout_factor_changed or posedge _check_t0_values )
    begin
        if (config_burst_timeout_factor_changed == 1'b1)
        begin
            axi_get_config_burst_timeout_factor_into_SystemVerilog( _interface_ref, config_burst_timeout_factor ); // DPI call to imported task
            config_burst_timeout_factor_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_AWVALID_assertion_to_AWREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_AWVALID_assertion_to_AWREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_AWVALID_assertion_to_AWREADY_into_SystemVerilog( _interface_ref, config_max_latency_AWVALID_assertion_to_AWREADY ); // DPI call to imported task
            config_max_latency_AWVALID_assertion_to_AWREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_ARVALID_assertion_to_ARREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_ARVALID_assertion_to_ARREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_ARVALID_assertion_to_ARREADY_into_SystemVerilog( _interface_ref, config_max_latency_ARVALID_assertion_to_ARREADY ); // DPI call to imported task
            config_max_latency_ARVALID_assertion_to_ARREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_RVALID_assertion_to_RREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_RVALID_assertion_to_RREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_RVALID_assertion_to_RREADY_into_SystemVerilog( _interface_ref, config_max_latency_RVALID_assertion_to_RREADY ); // DPI call to imported task
            config_max_latency_RVALID_assertion_to_RREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_BVALID_assertion_to_BREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_BVALID_assertion_to_BREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_BVALID_assertion_to_BREADY_into_SystemVerilog( _interface_ref, config_max_latency_BVALID_assertion_to_BREADY ); // DPI call to imported task
            config_max_latency_BVALID_assertion_to_BREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_WVALID_assertion_to_WREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_WVALID_assertion_to_WREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_WVALID_assertion_to_WREADY_into_SystemVerilog( _interface_ref, config_max_latency_WVALID_assertion_to_WREADY ); // DPI call to imported task
            config_max_latency_WVALID_assertion_to_WREADY_changed = 1'b0;
        end
    end

    always @(posedge config_master_error_position_changed or posedge _check_t0_values )
    begin
        if (config_master_error_position_changed == 1'b1)
        begin
            axi_get_config_master_error_position_into_SystemVerilog( _interface_ref, config_master_error_position ); // DPI call to imported task
            config_master_error_position_changed = 1'b0;
        end
    end

    always @(posedge config_setup_time_changed or posedge _check_t0_values )
    begin
        if (config_setup_time_changed == 1'b1)
        begin
            axi_get_config_setup_time_into_SystemVerilog( _interface_ref, config_setup_time ); // DPI call to imported task
            config_setup_time_changed = 1'b0;
        end
    end

    always @(posedge config_hold_time_changed or posedge _check_t0_values )
    begin
        if (config_hold_time_changed == 1'b1)
        begin
            axi_get_config_hold_time_into_SystemVerilog( _interface_ref, config_hold_time ); // DPI call to imported task
            config_hold_time_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_wr_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_wr_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_wr_into_SystemVerilog( _interface_ref, config_max_outstanding_wr ); // DPI call to imported task
            config_max_outstanding_wr_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_rd_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_rd_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_rd_into_SystemVerilog( _interface_ref, config_max_outstanding_rd ); // DPI call to imported task
            config_max_outstanding_rd_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_rw_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_rw_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_rw_into_SystemVerilog( _interface_ref, config_max_outstanding_rw ); // DPI call to imported task
            config_max_outstanding_rw_changed = 1'b0;
        end
    end

    always @(posedge config_is_issuing_changed or posedge _check_t0_values )
    begin
        if (config_is_issuing_changed == 1'b1)
        begin
            axi_get_config_is_issuing_into_SystemVerilog( _interface_ref, config_is_issuing ); // DPI call to imported task
            config_is_issuing_changed = 1'b0;
        end
    end


// Timeless transaction interface support

    // assocative array of event indexed by unique_id(int)
    event assoc_timeless_comm_array[int];

    // these three functions are used by the timeless_trans_control event loop:
    // 1. initialise the loop
    import "DPI-C" context axi_start_next_timeless_trans = function void axi_start_next_timeless_trans();
    // 2. get next completed timeless transaction, returns null at the end
    import "DPI-C" context axi_get_next_timeless_trans = function int axi_get_next_timeless_trans();
    // 3. reset loop and empty the list
    import "DPI-C" context axi_end_next_timeless_trans = function void axi_end_next_timeless_trans();
    // could do above a little more efficiently by having each 'get' also remove the element so won't need an 'end'?

    // when timeless transaction monitor goes to 1 ..... trigger all the events associated with each transaction
    always @(posedge timeless_trans_control)
    begin
        int _trans_id ;
        // initialise C++ list
        axi_start_next_timeless_trans() ; 
        // loop round the list, triggering all associated events
        for ( _trans_id= axi_get_next_timeless_trans() ;
              _trans_id != 0 ;
              _trans_id= axi_get_next_timeless_trans() )
        begin
            if ( assoc_timeless_comm_array.exists( _trans_id ) )
            begin
                // trigger the event
                -> assoc_timeless_comm_array[_trans_id] ;
                // the _END_ deletes it from the array after checking existance ...
                // - that's two accesses to the array here and two in the END, there must be a more efficient way! (Could do it in C++)
            end
            else
            begin
                // survivable (?) error - a non-null handle returned which isn't in the array!
                $display("Transaction WARNING @ %t: %m - unknown unique_id received from Adaptor.",$time);
            end
        end
        // completed C++ list
        axi_end_next_timeless_trans() ; 
        timeless_trans_control= 0 ;
    end

    //--------------------------------------------------------------------------------
    // Task which blocks and outputs an error if the interface has not initialized properly
    //--------------------------------------------------------------------------------

    task _initialized();
        if (_interface_ref == 0)
        begin
            $display("Error: %m - Questa Verification IP failed to initialise. Please check questa_mvc.log for details");
            wait(_interface_ref!=0);
        end
    endtask

endinterface

`endif // MODEL_TECH
`ifdef INCA
// *****************************************************************************
//
// Copyright 2007-2016 Mentor Graphics Corporation
// All Rights Reserved.
//
// THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE PROPERTY OF
// MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS.
//
// *****************************************************************************
// SystemVerilog           Version: 20160107
// *****************************************************************************

import QUESTA_MVC::questa_mvc_reporter;
import QUESTA_MVC::questa_mvc_item_comms_semantic;
import QUESTA_MVC::questa_mvc_edge;
import QUESTA_MVC::QUESTA_MVC_POSEDGE;
import QUESTA_MVC::QUESTA_MVC_NEGEDGE;
import QUESTA_MVC::QUESTA_MVC_ANYEDGE;
import QUESTA_MVC::QUESTA_MVC_0_TO_1_EDGE;
import QUESTA_MVC::QUESTA_MVC_1_TO_0_EDGE;


(* cy_so="libaxi_IN_SystemVerilog_MTI_full" *)
(* on_lib_load="axi_IN_SystemVerilog_load" *)

interface mgc_common_axi #(int AXI_ADDRESS_WIDTH = 64, int AXI_RDATA_WIDTH = 1024, int AXI_WDATA_WIDTH = 1024, int AXI_ID_WIDTH = 18)
    (input wire iACLK, input wire iARESETn);

    //-------------------------------------------------------------------------
    //
    // Group: AXI Signals
    //
    //-------------------------------------------------------------------------



    //-------------------------------------------------------------------------
    // Private wires
    //-------------------------------------------------------------------------
    wire ACLK;
    wire ARESETn;
    wire AWVALID;
    wire [((AXI_ADDRESS_WIDTH) - 1):0]  AWADDR;
    wire [3:0] AWLEN;
    wire [2:0] AWSIZE;
    wire [1:0] AWBURST;
    wire [1:0] AWLOCK;
    wire [3:0] AWCACHE;
    wire [2:0] AWPROT;
    wire [((AXI_ID_WIDTH) - 1):0]  AWID;
    wire AWREADY;
    wire [7:0] AWUSER;
    wire ARVALID;
    wire [((AXI_ADDRESS_WIDTH) - 1):0]  ARADDR;
    wire [3:0] ARLEN;
    wire [2:0] ARSIZE;
    wire [1:0] ARBURST;
    wire [1:0] ARLOCK;
    wire [3:0] ARCACHE;
    wire [2:0] ARPROT;
    wire [((AXI_ID_WIDTH) - 1):0]  ARID;
    wire ARREADY;
    wire [7:0] ARUSER;
    wire RVALID;
    wire RLAST;
    wire [((AXI_RDATA_WIDTH) - 1):0]  RDATA;
    wire [1:0] RRESP;
    wire [((AXI_ID_WIDTH) - 1):0]  RID;
    wire RREADY;
    wire [7:0] RUSER;
    wire WVALID;
    wire WLAST;
    wire [((AXI_WDATA_WIDTH) - 1):0]  WDATA;
    wire [(((AXI_WDATA_WIDTH / 8)) - 1):0]  WSTRB;
    wire [((AXI_ID_WIDTH) - 1):0]  WID;
    wire WREADY;
    wire [7:0] WUSER;
    wire BVALID;
    wire [1:0] BRESP;
    wire [((AXI_ID_WIDTH) - 1):0]  BID;
    wire BREADY;
    wire [7:0] BUSER;



    // Propagate global signals onto interface wires
    assign ACLK = iACLK;
    assign ARESETn = iARESETn;

    // Variable: config_write_ctrl_to_data_mintime
    //
    // 
    // Sets the delay from start of address phase to start of data phase in a write 
    // transaction (in terms of ACLK).
    // 
    // Default: 1 
    // 
    // This configuration variable has been deprecated and is maintained 
    // for backward compatibility. However, you can use ~write_address_to_data_delay~ 
    // configuration variable to control the delay between a write address phase 
    // and a write data phase.
    // 
    //
    int unsigned config_write_ctrl_to_data_mintime;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Enables
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_enable_all_assertions
    //
    // 
    // Enables all protocol assertions. 
    // 
    // Default: 1
    // 
    //
    // mentor configurator specification name "Enable all protocol assertions"
    bit config_enable_all_assertions;

    // Variable: config_enable_assertion
    //
    // 
    // Enables individual protocol assertion.
    // This variable controls whether specific assertion within QVIP (of type <axi_assertion_e>) is enabled or disabled.
    // Individual assertion can be disabled as follows:-
    // //-----------------------------------------------------------------------
    // // < BFM interface>.set_config_enable_assertion_index1(<name of assertion>,1'b0);
    // //-----------------------------------------------------------------------
    // 
    // For example, the assertion AXI_READ_DATA_UNKN is disabled as follows:
    // <bfm>.set_config_enable_assertion_index1(AXI_READ_DATA_UNKN, 1'b0); 
    // 
    // Here bfm is the AXI interface instance name for which the assertion to be disabled. 
    // 
    // Default: All assertions are enabled
    //   
    // 
    //
    // mentor configurator specification name "Enable individual protocol assertion"
    bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Slave behavior control
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_support_exclusive_access
    //
    // 
    // Enables exclusive transactions support for slave.
    // If disabled, every exclusive read/write returns an OKAY response,
    // and exclusive write updates memory. 
    // 
    // Default: 1  
    // 
    //
    // mentor configurator specification name "Enable exclusive transaction support"
    bit config_support_exclusive_access;

    // Variable: config_read_data_reordering_depth
    //
    // 
    // Sets the maximum number of different read transaction addresses for which read 
    // data(response) can be sent in any order from slave. 
    // 
    // Default: 2 ** AXI_ID_WIDTH
    // 
    //
    // mentor configurator specification name "Read data reordering depth"
    int unsigned config_read_data_reordering_depth;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Timeout control
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_max_transaction_time_factor
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) for any complete read or write transaction, which
    // includes time period for all individual phases of transaction. 
    // 
    // Default: 100000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout for complete read/write transaction"
    int unsigned config_max_transaction_time_factor;

    // Variable: config_timeout_max_data_transfer
    //
    //  
    // Sets maximum number of write data beats in a write data burst. 
    // 
    // Default: 1024  
    // 
    //
    // mentor configurator specification name "Maximum number of data beats in a write data burst"
    int config_timeout_max_data_transfer;

    // Variable: config_burst_timeout_factor
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) between individual phases of a transaction. 
    // 
    // Default: 10000 clock cycles 
    // 
    //
    // mentor configurator specification name "Burst timeout between individual phases of a transaction"
    int unsigned config_burst_timeout_factor;

    // Variable: config_max_latency_AWVALID_assertion_to_AWREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of AWVALID to assertion of AWREADY.
    // An error message AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID is generated if AWREADY is not asserted
    // after assertion of AWVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from AWVALID to AWREADY assertion"
    int unsigned config_max_latency_AWVALID_assertion_to_AWREADY;

    // Variable: config_max_latency_ARVALID_assertion_to_ARREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of ARVALID to assertion of ARREADY.
    // An error message AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID is generated if ARREADY is not asserted
    // after assertion of ARVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from ARVALID to ARREADY assertion"
    int unsigned config_max_latency_ARVALID_assertion_to_ARREADY;

    // Variable: config_max_latency_RVALID_assertion_to_RREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of RVALID to assertion of RREADY.
    // An error message AXI_RREADY_NOT_ASSERTED_AFTER_RVALID is generated if RREADY is not asserted
    // after assertion of RVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from RVALID to RREADY assertion"
    int unsigned config_max_latency_RVALID_assertion_to_RREADY;

    // Variable: config_max_latency_BVALID_assertion_to_BREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of BVALID to assertion of BREADY.
    // An error message AXI_BREADY_NOT_ASSERTED_AFTER_BVALID is generated if BREADY is not asserted
    // after assertion of BVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from BVALID to BREADY assertion"
    int unsigned config_max_latency_BVALID_assertion_to_BREADY;

    // Variable: config_max_latency_WVALID_assertion_to_WREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of WVALID to assertion of WREADY.
    // An error message AXI_WREADY_NOT_ASSERTED_AFTER_WVALID is generated if WREADY is not asserted
    // after assertion of WVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from WVALID to WREADY assertion"
    int unsigned config_max_latency_WVALID_assertion_to_WREADY;

    // Variable: config_setup_time
    //
    // 
    // Sets number of simulation time units from the setup time to the active 
    // clock edge of ACLK. The setup time will always be less than the time period
    // of the clock. 
    // 
    // Default: 0
    // 
    //
    // Note - This configuration variable is used in an expression involving time precision.
    //        To ensure its value is correct, use questa_mvc_sv_convert_to_precision API of QUESTA_MVC package.
    //
    int config_setup_time;

    // Variable: config_hold_time
    //
    // 
    // Sets number of simulation time units from the hold time to the active 
    // clock edge of ACLK. 
    // 
    // Default: 0
    // 
    //
    // Note - This configuration variable is used in an expression involving time precision.
    //        To ensure its value is correct, use questa_mvc_sv_convert_to_precision API of QUESTA_MVC package.
    //
    int config_hold_time;

    // Variable: config_max_outstanding_wr
    //
    // Configures maximum possible outstanding Write transactions
    //
    int config_max_outstanding_wr;

    // Variable: config_max_outstanding_rd
    //
    // Configures maximum possible outstanding Read transactions
    //
    int config_max_outstanding_rd;

    // Variable: config_max_outstanding_rw
    //
    // Configures maximum possible outstanding Combined (Read and Write) transactions
    //
    int config_max_outstanding_rw;

    // Variable: config_is_issuing
    //
    // Enables Master component to use "config_max_outstanding_wr/config_max_outstanding_rd/config_max_outstanding_rw" variables for transaction issuing capability when set to true
    //
    bit config_is_issuing;


    //-------------------------------------------------------------------------
    // Deprecated variables - writing to these variables will cause a warning to be issued.
    //-------------------------------------------------------------------------
    bit config_master_write_delay;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr;
    axi_error_e config_master_error_position;
    //------------------------------------------------------------------------------
    // Group:- Interface ends
    //------------------------------------------------------------------------------
    //
    longint axi_master_end;


    // Function:- get_axi_master_end
    //
    // Returns a handle to the <master> end of this instance of the <axi> interface.

    function longint get_axi_master_end();
        return axi_master_end;
    endfunction

    longint axi_slave_end;


    // Function:- get_axi_slave_end
    //
    // Returns a handle to the <slave> end of this instance of the <axi> interface.

    function longint get_axi_slave_end();
        return axi_slave_end;
    endfunction

    longint axi_clock_source_end;


    // Function:- get_axi_clock_source_end
    //
    // Returns a handle to the <clock_source> end of this instance of the <axi> interface.

    function longint get_axi_clock_source_end();
        return axi_clock_source_end;
    endfunction

    longint axi_reset_source_end;


    // Function:- get_axi_reset_source_end
    //
    // Returns a handle to the <reset_source> end of this instance of the <axi> interface.

    function longint get_axi_reset_source_end();
        return axi_reset_source_end;
    endfunction

    longint axi__monitor_end;


    // Function:- get_axi__monitor_end
    //
    // Returns a handle to the <_monitor> end of this instance of the <axi> interface.

    function longint get_axi__monitor_end();
        return axi__monitor_end;
    endfunction


    // Group:- Abstraction Levels
    // 
    // These functions are used set or get the abstraction levels of an interface end.
    // See <Abstraction Levels of Interface Ends> for more details on the meaning of
    // TLM or WLM connected and the valid combinations.


    //-------------------------------------------------------------------------
    // Function:- axi_set_master_abstraction_level
    //
    //     Function to set whether the <master> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_master_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_master_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_master_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <master> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_master_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_master_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_slave_abstraction_level
    //
    //     Function to set whether the <slave> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_slave_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_slave_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_slave_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <slave> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_slave_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_slave_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_clock_source_abstraction_level
    //
    //     Function to set whether the <clock_source> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_clock_source_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_clock_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_clock_source_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <clock_source> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_clock_source_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_clock_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_reset_source_abstraction_level
    //
    //     Function to set whether the <reset_source> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_reset_source_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_reset_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_reset_source_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <reset_source> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_reset_source_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_reset_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    import "DPI-C" context function longint axi_initialise_SystemVerilog
    (
        int    usage_code,
        string iface_version,
        output longint master_end,
        output longint slave_end,
        output longint clock_source_end,
        output longint reset_source_end,
        output longint _monitor_end,
        input int AXI_ADDRESS_WIDTH,
        input int AXI_RDATA_WIDTH,
        input int AXI_WDATA_WIDTH,
        input int AXI_ID_WIDTH
    );

    `ifndef MVC_axi_VERSION
    `define MVC_axi_VERSION ""
    `endif
    // Handle to the linkage
    (* elab_init *) longint _interface_ref =
                                axi_initialise_SystemVerilog
                                (
                                    18102076,
                                    `MVC_axi_VERSION,
                                    axi_master_end,
                                    axi_slave_end,
                                    axi_clock_source_end,
                                    axi_reset_source_end,
                                    axi__monitor_end,
                                    AXI_ADDRESS_WIDTH,
                                    AXI_RDATA_WIDTH,
                                    AXI_WDATA_WIDTH,
                                    AXI_ID_WIDTH
                                ); // DPI call to create transactor (called at
                                     // elaboration time as initialiser)

        bit report_available;

        // Function for getting a message from QUESTA_MVC. Returns 1 if a message was returned, 0 otherwise.
        import "DPI-C" questa_mvc_sv_get_report =  function bit get_report( input longint iface_ref,input longint recipient,
                                     output string category,     output string objectName,
                                     output string instanceName, output string error_no,
                                     output string typ,          output string mess );
        questa_mvc_reporter endPoint[longint];
        initial report_available = 0;

        always @report_available
        begin
            longint recipient;
            string category;
            string objectName;
            string instanceName;
            string severity;
            string mess;
            string error_no;

            if ( endPoint.first( recipient ) )
              begin
                do
                  begin
                      while ( get_report( _interface_ref, recipient, category, objectName, instanceName, error_no, severity, mess ) )
                        begin
                          endPoint[recipient].report_message( category, "axi", 0, objectName, instanceName, error_no, severity, mess );
                        end
                  end
                while (endPoint.next(recipient));
              end
            report_available = 0;
        end

        import "DPI-C" context questa_mvc_register_end_point = function void questa_mvc_register_end_point( input longint iface_ref, input longint as_end, input string name );

        // A function for registering a reporter to capture any reports coming from as_end
        function automatic void register_end_point( input longint as_end, input questa_mvc_reporter rep = null );
            if ( rep != null )
              begin
                if ( ( rep.name == "" ) || ( rep.name == "NULL" ) )
                  begin
                    $display("Error: %m: Reporter passed to register_end_point has a reserved name. Neither an empty string nor the string 'NULL' can be used.");
                  end
                else
                  begin
                    questa_mvc_register_end_point( _interface_ref, as_end, rep.name );
                    endPoint[as_end] = rep;
                  end
              end
            else
              begin
                questa_mvc_register_end_point( _interface_ref, as_end, "NULL" );
                endPoint.delete( as_end );
              end
        endfunction

    //-------------------------------------------------------------------------
    //
    // Group:- Registering Reports
    //
    //
    // The following methods are used to register a custom reporting object as
    // described in the MVC base library section, <Customizing Error-Reporting>.
    // 
    //-------------------------------------------------------------------------

    function void register_interface_reporter( input questa_mvc_reporter _rep = null );
        register_end_point( _interface_ref, _rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_master_reporter
    //
    // Function used to register a reporter for the <master> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the master end.
    //
    function void register_master_reporter
    (
        input questa_mvc_reporter rep = null
    );
        register_end_point( axi_master_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_slave_reporter
    //
    // Function used to register a reporter for the <slave> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the slave end.
    //
    function void register_slave_reporter
    (
        input questa_mvc_reporter rep = null
    );
        register_end_point( axi_slave_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_clock_source_reporter
    //
    // Function used to register a reporter for the <clock_source> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the clock_source end.
    //
    function void register_clock_source_reporter
    (
        input questa_mvc_reporter rep = null
    );
        register_end_point( axi_clock_source_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_reset_source_reporter
    //
    // Function used to register a reporter for the <reset_source> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the reset_source end.
    //
    function void register_reset_source_reporter
    (
        input questa_mvc_reporter rep = null
    );
        register_end_point( axi_reset_source_end, rep );
    endfunction


    //-------------------------------------------------------------------------
    //
    // Group:- BFM Utility/Convenience Methods
    //
    // This is the group of utility functions provided by the QVIP BFM to
    // communicate from the SV world to the QVIP BFM.
    // This set of APIs can be used to either get status/statistics
    // information from the BFM or to set values in a particular database 
    // in the BFM. Please refer to individual functions for more information.
    //
    //-------------------------------------------------------------------------

    export "DPI-C" axi_get_temp_static_fn_rd_txn_valid_lanes_valid_lanes = function axi_get_temp_static_fn_rd_txn_valid_lanes_valid_lanes;
    export "DPI-C" axi_set_temp_static_fn_rd_txn_valid_lanes_valid_lanes = function axi_set_temp_static_fn_rd_txn_valid_lanes_valid_lanes;
    bit [((AXI_RDATA_WIDTH / 8) - 1):0] temp_static_fn_rd_txn_valid_lanes_valid_lanes [];
    function void axi_get_temp_static_fn_rd_txn_valid_lanes_valid_lanes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_fn_rd_txn_valid_lanes_valid_lanes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_fn_rd_txn_valid_lanes_valid_lanes( input int _d1, input int _d2, input bit _value );
        temp_static_fn_rd_txn_valid_lanes_valid_lanes[_d1][_d2] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_rd_txn_valid_lanes
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get valid strobes/lanes value for each of the read data beat
    //     at end of read transaction.
    // 
    //     Please note that this function should be called after completion of a read
    //     transaction.
    // 
    //     Output of the function:
    //     valid_lanes - Valid strobes value for each read data beat
    //    
    function automatic void fn_rd_txn_valid_lanes
    (
        ref bit [((AXI_RDATA_WIDTH / 8) - 1):0] valid_lanes []
    );
        temp_static_fn_rd_txn_valid_lanes_valid_lanes = new[valid_lanes.size()];
         fn_rd_txn_valid_lanes_C();
        valid_lanes = temp_static_fn_rd_txn_valid_lanes_valid_lanes;
    endfunction

    export "DPI-C" axi_get_temp_static_fn_get_wdata_phase_info_id = function axi_get_temp_static_fn_get_wdata_phase_info_id;
    export "DPI-C" axi_set_temp_static_fn_get_wdata_phase_info_id = function axi_set_temp_static_fn_get_wdata_phase_info_id;
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_fn_get_wdata_phase_info_id;
    function void axi_get_temp_static_fn_get_wdata_phase_info_id( input int _d1, output bit  _value );
        _value = temp_static_fn_get_wdata_phase_info_id[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_wdata_phase_info_id( input int _d1, input bit  _value );
        temp_static_fn_get_wdata_phase_info_id[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_get_wdata_phase_info_beat_addr = function axi_get_temp_static_fn_get_wdata_phase_info_beat_addr;
    export "DPI-C" axi_set_temp_static_fn_get_wdata_phase_info_beat_addr = function axi_set_temp_static_fn_get_wdata_phase_info_beat_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_get_wdata_phase_info_beat_addr;
    function void axi_get_temp_static_fn_get_wdata_phase_info_beat_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_get_wdata_phase_info_beat_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_wdata_phase_info_beat_addr( input int _d1, input bit  _value );
        temp_static_fn_get_wdata_phase_info_beat_addr[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_get_wdata_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get information corresponding to a write data beat.
    // 
    //     Input:
    //     id         - ID of the write data beat
    //     wdata_last - assigned to ~last~ attribute of the write data beat
    // 
    //     Output:
    //     waddr_rcvd   - Indicates if corresponding write address phase is received
    //     burst_length - Burst length attribute of the corresponding address phase
    //     beat_num     - Write data beat number of the corresponding write data burst
    //     beat_addr    - Corresponding beat address
    // 
    //     Please note that this function should be called at the completion of write
    //     data beat.
    //    
    function automatic void fn_get_wdata_phase_info
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit wdata_last,
        inout bit waddr_rcvd,
        output bit [3:0] burst_length,
        output int beat_num,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  beat_addr
    );
        temp_static_fn_get_wdata_phase_info_id = id;
         fn_get_wdata_phase_info_C(wdata_last,waddr_rcvd,burst_length,beat_num);
        beat_addr = temp_static_fn_get_wdata_phase_info_beat_addr;
    endfunction

    export "DPI-C" axi_get_temp_static_fn_get_wresp_phase_info_wresp_corr_addr = function axi_get_temp_static_fn_get_wresp_phase_info_wresp_corr_addr;
    export "DPI-C" axi_set_temp_static_fn_get_wresp_phase_info_wresp_corr_addr = function axi_set_temp_static_fn_get_wresp_phase_info_wresp_corr_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_get_wresp_phase_info_wresp_corr_addr;
    function void axi_get_temp_static_fn_get_wresp_phase_info_wresp_corr_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_get_wresp_phase_info_wresp_corr_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_wresp_phase_info_wresp_corr_addr( input int _d1, input bit  _value );
        temp_static_fn_get_wresp_phase_info_wresp_corr_addr[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_get_wresp_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get address attribute of write address phase corresponding
    //     to write response phase that just completed.
    // 
    //     Please note that this function should be called after completion of a write
    //     response phase.
    // 
    //     Output of the function:
    //     wresp_corr_addr - ~addr~ attribute of the address phase corresponding to
    //                       this write response phase
    //    
    function automatic void fn_get_wresp_phase_info
    (
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  wresp_corr_addr
    );
         fn_get_wresp_phase_info_C();
        wresp_corr_addr = temp_static_fn_get_wresp_phase_info_wresp_corr_addr;
    endfunction

    export "DPI-C" axi_get_temp_static_fn_get_rdata_phase_info_id = function axi_get_temp_static_fn_get_rdata_phase_info_id;
    export "DPI-C" axi_set_temp_static_fn_get_rdata_phase_info_id = function axi_set_temp_static_fn_get_rdata_phase_info_id;
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_fn_get_rdata_phase_info_id;
    function void axi_get_temp_static_fn_get_rdata_phase_info_id( input int _d1, output bit  _value );
        _value = temp_static_fn_get_rdata_phase_info_id[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_rdata_phase_info_id( input int _d1, input bit  _value );
        temp_static_fn_get_rdata_phase_info_id[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_get_rdata_phase_info_beat_strobes = function axi_get_temp_static_fn_get_rdata_phase_info_beat_strobes;
    export "DPI-C" axi_set_temp_static_fn_get_rdata_phase_info_beat_strobes = function axi_set_temp_static_fn_get_rdata_phase_info_beat_strobes;
    bit [((AXI_RDATA_WIDTH / 8) - 1):0]  temp_static_fn_get_rdata_phase_info_beat_strobes;
    function void axi_get_temp_static_fn_get_rdata_phase_info_beat_strobes( input int _d1, output bit  _value );
        _value = temp_static_fn_get_rdata_phase_info_beat_strobes[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_rdata_phase_info_beat_strobes( input int _d1, input bit  _value );
        temp_static_fn_get_rdata_phase_info_beat_strobes[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_get_rdata_phase_info_beat_addr = function axi_get_temp_static_fn_get_rdata_phase_info_beat_addr;
    export "DPI-C" axi_set_temp_static_fn_get_rdata_phase_info_beat_addr = function axi_set_temp_static_fn_get_rdata_phase_info_beat_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_get_rdata_phase_info_beat_addr;
    function void axi_get_temp_static_fn_get_rdata_phase_info_beat_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_get_rdata_phase_info_beat_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_rdata_phase_info_beat_addr( input int _d1, input bit  _value );
        temp_static_fn_get_rdata_phase_info_beat_addr[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_get_rdata_phase_info_txn_addr = function axi_get_temp_static_fn_get_rdata_phase_info_txn_addr;
    export "DPI-C" axi_set_temp_static_fn_get_rdata_phase_info_txn_addr = function axi_set_temp_static_fn_get_rdata_phase_info_txn_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_get_rdata_phase_info_txn_addr;
    function void axi_get_temp_static_fn_get_rdata_phase_info_txn_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_get_rdata_phase_info_txn_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_rdata_phase_info_txn_addr( input int _d1, input bit  _value );
        temp_static_fn_get_rdata_phase_info_txn_addr[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_get_rdata_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get information corresponding to a read data beat.
    // 
    //     Input:
    //     id         - ID of the read data beat
    // 
    //     Output:
    //     burst_length - Burst length attribute of the corresponding read address phase
    //     beat_num     - Read data beat number of the corresponding read data burst
    //     beat_strobes - Valid lanes in the read data beat
    //     beat_addr    - Corresponding beat address
    // 
    //     Please note that this function should be called at the completion of read
    //     data beat.
    //    
    function automatic void fn_get_rdata_phase_info
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit rdata_last,
        output bit [3:0] burst_length,
        output int beat_num,
        output bit [((AXI_RDATA_WIDTH / 8) - 1):0]  beat_strobes,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  beat_addr,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  txn_addr
    );
        temp_static_fn_get_rdata_phase_info_id = id;
         fn_get_rdata_phase_info_C(rdata_last,burst_length,beat_num);
        beat_strobes = temp_static_fn_get_rdata_phase_info_beat_strobes;
        beat_addr = temp_static_fn_get_rdata_phase_info_beat_addr;
        txn_addr = temp_static_fn_get_rdata_phase_info_txn_addr;
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_get_max_os_per_id
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function gets the maximum number of outstanding write phases of a particular ID
    // from among all AWID, WID values.
    //  
    // Inputs:
    // max_waddr_os - The maximum number of address phases outstanding from among all AWID
    // max_wdata_os - The maximum number of data bursts outstanding from among all WID
    // 
    // For example, 5 write address phases are outstanding with ID 3, and 
    // 7 write address phases are outstanding with ID 2. No other address phase is there
    // and 0 write data phases are received.
    // 
    // The return values would be such that:
    // max_waddr_os = 7
    // max_wdata_os = 0
    // 
    function automatic void fn_get_max_os_per_id
    (
        output int max_waddr_os,
        output int max_wdata_os
    );
         fn_get_max_os_per_id_C(max_waddr_os,max_wdata_os);
    endfunction

    export "DPI-C" axi_get_temp_static_get_rw_txns_in_prog_id = function axi_get_temp_static_get_rw_txns_in_prog_id;
    export "DPI-C" axi_set_temp_static_get_rw_txns_in_prog_id = function axi_set_temp_static_get_rw_txns_in_prog_id;
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_get_rw_txns_in_prog_id;
    function void axi_get_temp_static_get_rw_txns_in_prog_id( input int _d1, output bit  _value );
        _value = temp_static_get_rw_txns_in_prog_id[_d1];
    endfunction
    function void axi_set_temp_static_get_rw_txns_in_prog_id( input int _d1, input bit  _value );
        temp_static_get_rw_txns_in_prog_id[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: get_rw_txns_in_prog
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function gets the number of various outstanding transactions at a time.
    // 
    // Inputs:
    // id  - The AWID/ARID/WID of the transaction whose details are required.
    // txn_counts - The statistics of the number of outstanding transactions
    function automatic void get_rw_txns_in_prog
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_rw_txn_counts_s txn_counts
    );
        temp_static_get_rw_txns_in_prog_id = id;
         get_rw_txns_in_prog_C(txn_counts);
    endfunction

    export "DPI-C" axi_get_temp_static_fn_add_addr_map_entry_addr = function axi_get_temp_static_fn_add_addr_map_entry_addr;
    export "DPI-C" axi_set_temp_static_fn_add_addr_map_entry_addr = function axi_set_temp_static_fn_add_addr_map_entry_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_add_addr_map_entry_addr;
    function void axi_get_temp_static_fn_add_addr_map_entry_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_add_addr_map_entry_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_add_addr_map_entry_addr( input int _d1, input bit  _value );
        temp_static_fn_add_addr_map_entry_addr[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_add_addr_map_entry
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets address map fields inside internal BFM. 
    // 
    // Inputs:
    // region - Region name 
    // addr - Start address of region
    // size - Size of address region
    function automatic void fn_add_addr_map_entry
    (
        input string region,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input longint unsigned size
    );
        temp_static_fn_add_addr_map_entry_addr = addr;
         fn_add_addr_map_entry_C(region,size);
    endfunction

    export "DPI-C" axi_get_temp_static_fn_add_wr_delay_data2data = function axi_get_temp_static_fn_add_wr_delay_data2data;
    export "DPI-C" axi_set_temp_static_fn_add_wr_delay_data2data = function axi_set_temp_static_fn_add_wr_delay_data2data;
    int unsigned temp_static_fn_add_wr_delay_data2data[];
    function void axi_get_temp_static_fn_add_wr_delay_data2data( input int _d1, output int unsigned _value );
        _value = temp_static_fn_add_wr_delay_data2data[_d1];
    endfunction
    function void axi_set_temp_static_fn_add_wr_delay_data2data( input int _d1, input int unsigned _value );
        temp_static_fn_add_wr_delay_data2data[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_add_wr_delay
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets delay values for write address-data pair and 
    // between write data beats, initiated by master end. 
    // 
    // Inputs:
    // region - Region value for which write delays are to be inserted
    // id - Write transaction's id (AWID) for which delays are to be inserted
    // addr2data - Delays to be inserted between write address and data phase.
    // data2data - Delays to be inserted between data beats
    function automatic void fn_add_wr_delay
    (
        input string region,
        input bit [17:0] id,
        input int unsigned addr2data,
        ref int unsigned data2data[]
    );
        int tmp_data2data_DIMS0;
        tmp_data2data_DIMS0 = data2data.size();
        temp_static_fn_add_wr_delay_data2data = data2data;
         fn_add_wr_delay_C(region,id,addr2data,tmp_data2data_DIMS0);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_delete_wr_delay
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function deletes delay values for a region-id pair
    // 
    // Inputs:
    // region - Region value for which write delays are to be inserted
    // id - Write transaction's id (AWID) for which delays are to be inserted
    // addr2data - Delays to be inserted between write address and data phase.
    // data2data - Delays to be inserted between data beats
    function automatic void fn_delete_wr_delay
    (
        input string region,
        input bit [17:0] id
    );
         fn_delete_wr_delay_C(region,id);
    endfunction

    export "DPI-C" axi_get_temp_static_fn_set_wr_def_delays_min_data2data = function axi_get_temp_static_fn_set_wr_def_delays_min_data2data;
    export "DPI-C" axi_set_temp_static_fn_set_wr_def_delays_min_data2data = function axi_set_temp_static_fn_set_wr_def_delays_min_data2data;
    int unsigned temp_static_fn_set_wr_def_delays_min_data2data[];
    function void axi_get_temp_static_fn_set_wr_def_delays_min_data2data( input int _d1, output int unsigned _value );
        _value = temp_static_fn_set_wr_def_delays_min_data2data[_d1];
    endfunction
    function void axi_set_temp_static_fn_set_wr_def_delays_min_data2data( input int _d1, input int unsigned _value );
        temp_static_fn_set_wr_def_delays_min_data2data[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_set_wr_def_delays_max_data2data = function axi_get_temp_static_fn_set_wr_def_delays_max_data2data;
    export "DPI-C" axi_set_temp_static_fn_set_wr_def_delays_max_data2data = function axi_set_temp_static_fn_set_wr_def_delays_max_data2data;
    int unsigned temp_static_fn_set_wr_def_delays_max_data2data[];
    function void axi_get_temp_static_fn_set_wr_def_delays_max_data2data( input int _d1, output int unsigned _value );
        _value = temp_static_fn_set_wr_def_delays_max_data2data[_d1];
    endfunction
    function void axi_set_temp_static_fn_set_wr_def_delays_max_data2data( input int _d1, input int unsigned _value );
        temp_static_fn_set_wr_def_delays_max_data2data[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_set_wr_def_delays
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets default delay values for write address-data pair and data beats 
    // initiated by master end between input max. and min. values. In case non-randomized 
    // default value is desired, user can set max. and min. to same value.
    // 
    // Inputs:
    // min_addr2data - Minimum value of default delays to be inserted between write address and data phase.
    // min_data2data - Minimum value of default delays to be inserted between data beats
    // max_addr2data - Maximum value of default delays to be inserted between write address and data phase.
    // max_data2data - Maximum value of default delays to be inserted between data beats
    function automatic void fn_set_wr_def_delays
    (
        input int unsigned min_addr2data,
        ref int unsigned min_data2data[],
        input int unsigned max_addr2data,
        ref int unsigned max_data2data[]
    );
        int tmp_min_data2data_DIMS0;
        int tmp_max_data2data_DIMS0;
        tmp_min_data2data_DIMS0 = min_data2data.size();
        tmp_max_data2data_DIMS0 = max_data2data.size();
        temp_static_fn_set_wr_def_delays_min_data2data = min_data2data;
        temp_static_fn_set_wr_def_delays_max_data2data = max_data2data;
         fn_set_wr_def_delays_C(min_addr2data,tmp_min_data2data_DIMS0,max_addr2data,tmp_max_data2data_DIMS0);
    endfunction

    // Declare user visible wires variables, for non-continuous assignments.
    logic m_ACLK = 'z;
    logic m_ARESETn = 'z;
    logic m_AWVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  m_AWADDR = 'z;
    logic [3:0] m_AWLEN = 'z;
    logic [2:0] m_AWSIZE = 'z;
    logic [1:0] m_AWBURST = 'z;
    logic [1:0] m_AWLOCK = 'z;
    logic [3:0] m_AWCACHE = 'z;
    logic [2:0] m_AWPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_AWID = 'z;
    logic m_AWREADY = 'z;
    logic [7:0] m_AWUSER = 'z;
    logic m_ARVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  m_ARADDR = 'z;
    logic [3:0] m_ARLEN = 'z;
    logic [2:0] m_ARSIZE = 'z;
    logic [1:0] m_ARBURST = 'z;
    logic [1:0] m_ARLOCK = 'z;
    logic [3:0] m_ARCACHE = 'z;
    logic [2:0] m_ARPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_ARID = 'z;
    logic m_ARREADY = 'z;
    logic [7:0] m_ARUSER = 'z;
    logic m_RVALID = 'z;
    logic m_RLAST = 'z;
    logic [((AXI_RDATA_WIDTH) - 1):0]  m_RDATA = 'z;
    logic [1:0] m_RRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_RID = 'z;
    logic m_RREADY = 'z;
    logic [7:0] m_RUSER = 'z;
    logic m_WVALID = 'z;
    logic m_WLAST = 'z;
    logic [((AXI_WDATA_WIDTH) - 1):0]  m_WDATA = 'z;
    logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  m_WSTRB = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_WID = 'z;
    logic m_WREADY = 'z;
    logic [7:0] m_WUSER = 'z;
    logic m_BVALID = 'z;
    logic [1:0] m_BRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_BID = 'z;
    logic m_BREADY = 'z;
    logic [7:0] m_BUSER = 'z;

    // Forces a sweep through the wire change checkers at time 0 to get around
    // process kick-off order unknowns
    bit _check_t0_values;
    always_comb _check_t0_values = 1;

    // handle control
    longint last_handle = 0;

    longint last_start_time = 0;

    longint last_end_time = 0;

    export "DPI-C" axi_set_last_handle_and_times = function set_last_handle_and_times;

    function void set_last_handle_and_times(longint _handle, longint _start, longint _end);
        last_handle = _handle;
        last_start_time = _start;
        last_end_time = _end;
    endfunction


    function longint get_last_handle();
        return last_handle;
    endfunction


    function longint get_last_start_time();
        return last_start_time;
    endfunction


    function longint get_last_end_time();
        return last_end_time;
    endfunction


    //-------------------------------------------------------------------------
    // Tasks to wait for a number of specified edges on a wire
    //-------------------------------------------------------------------------


    //------------------------------------------------------------------------------
    // Function:- wait_for_ACLK
    //     Wait for the specified change on wire <axi::ACLK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ACLK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ACLK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ACLK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ACLK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ACLK === 0 );
                    @( ACLK );
                end
                while ( ACLK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ACLK === 1 );
                    @( ACLK );
                end
                while ( ACLK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARESETn
    //     Wait for the specified change on wire <axi::ARESETn>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARESETn( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARESETn);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARESETn);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARESETn);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARESETn === 0 );
                    @( ARESETn );
                end
                while ( ARESETn !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARESETn === 1 );
                    @( ARESETn );
                end
                while ( ARESETn !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWVALID
    //     Wait for the specified change on wire <axi::AWVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWVALID === 0 );
                    @( AWVALID );
                end
                while ( AWVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWVALID === 1 );
                    @( AWVALID );
                end
                while ( AWVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWADDR
    //     Wait for the specified change on wire <axi::AWADDR>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWADDR( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWADDR);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWADDR);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWADDR);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWADDR === 0 );
                    @( AWADDR );
                end
                while ( AWADDR !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWADDR === 1 );
                    @( AWADDR );
                end
                while ( AWADDR !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWADDR_index1
    //     Wait for the specified change on wire <axi::AWADDR>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWADDR_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWADDR[_this_dot_1] === 0 );
                    @( AWADDR[_this_dot_1] );
                end
                while ( AWADDR[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWADDR[_this_dot_1] === 1 );
                    @( AWADDR[_this_dot_1] );
                end
                while ( AWADDR[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLEN
    //     Wait for the specified change on wire <axi::AWLEN>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLEN( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLEN);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLEN);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLEN);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLEN === 0 );
                    @( AWLEN );
                end
                while ( AWLEN !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLEN === 1 );
                    @( AWLEN );
                end
                while ( AWLEN !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLEN_index1
    //     Wait for the specified change on wire <axi::AWLEN>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLEN_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLEN[_this_dot_1] === 0 );
                    @( AWLEN[_this_dot_1] );
                end
                while ( AWLEN[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLEN[_this_dot_1] === 1 );
                    @( AWLEN[_this_dot_1] );
                end
                while ( AWLEN[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWSIZE
    //     Wait for the specified change on wire <axi::AWSIZE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWSIZE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWSIZE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWSIZE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWSIZE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWSIZE === 0 );
                    @( AWSIZE );
                end
                while ( AWSIZE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWSIZE === 1 );
                    @( AWSIZE );
                end
                while ( AWSIZE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWSIZE_index1
    //     Wait for the specified change on wire <axi::AWSIZE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWSIZE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWSIZE[_this_dot_1] === 0 );
                    @( AWSIZE[_this_dot_1] );
                end
                while ( AWSIZE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWSIZE[_this_dot_1] === 1 );
                    @( AWSIZE[_this_dot_1] );
                end
                while ( AWSIZE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWBURST
    //     Wait for the specified change on wire <axi::AWBURST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWBURST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWBURST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWBURST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWBURST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWBURST === 0 );
                    @( AWBURST );
                end
                while ( AWBURST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWBURST === 1 );
                    @( AWBURST );
                end
                while ( AWBURST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWBURST_index1
    //     Wait for the specified change on wire <axi::AWBURST>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWBURST_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWBURST[_this_dot_1] === 0 );
                    @( AWBURST[_this_dot_1] );
                end
                while ( AWBURST[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWBURST[_this_dot_1] === 1 );
                    @( AWBURST[_this_dot_1] );
                end
                while ( AWBURST[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLOCK
    //     Wait for the specified change on wire <axi::AWLOCK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLOCK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLOCK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLOCK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLOCK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLOCK === 0 );
                    @( AWLOCK );
                end
                while ( AWLOCK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLOCK === 1 );
                    @( AWLOCK );
                end
                while ( AWLOCK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLOCK_index1
    //     Wait for the specified change on wire <axi::AWLOCK>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLOCK_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLOCK[_this_dot_1] === 0 );
                    @( AWLOCK[_this_dot_1] );
                end
                while ( AWLOCK[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLOCK[_this_dot_1] === 1 );
                    @( AWLOCK[_this_dot_1] );
                end
                while ( AWLOCK[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWCACHE
    //     Wait for the specified change on wire <axi::AWCACHE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWCACHE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWCACHE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWCACHE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWCACHE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWCACHE === 0 );
                    @( AWCACHE );
                end
                while ( AWCACHE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWCACHE === 1 );
                    @( AWCACHE );
                end
                while ( AWCACHE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWCACHE_index1
    //     Wait for the specified change on wire <axi::AWCACHE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWCACHE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWCACHE[_this_dot_1] === 0 );
                    @( AWCACHE[_this_dot_1] );
                end
                while ( AWCACHE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWCACHE[_this_dot_1] === 1 );
                    @( AWCACHE[_this_dot_1] );
                end
                while ( AWCACHE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWPROT
    //     Wait for the specified change on wire <axi::AWPROT>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWPROT( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWPROT);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWPROT);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWPROT);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWPROT === 0 );
                    @( AWPROT );
                end
                while ( AWPROT !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWPROT === 1 );
                    @( AWPROT );
                end
                while ( AWPROT !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWPROT_index1
    //     Wait for the specified change on wire <axi::AWPROT>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWPROT_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWPROT[_this_dot_1] === 0 );
                    @( AWPROT[_this_dot_1] );
                end
                while ( AWPROT[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWPROT[_this_dot_1] === 1 );
                    @( AWPROT[_this_dot_1] );
                end
                while ( AWPROT[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWID
    //     Wait for the specified change on wire <axi::AWID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWID === 0 );
                    @( AWID );
                end
                while ( AWID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWID === 1 );
                    @( AWID );
                end
                while ( AWID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWID_index1
    //     Wait for the specified change on wire <axi::AWID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWID[_this_dot_1] === 0 );
                    @( AWID[_this_dot_1] );
                end
                while ( AWID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWID[_this_dot_1] === 1 );
                    @( AWID[_this_dot_1] );
                end
                while ( AWID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWREADY
    //     Wait for the specified change on wire <axi::AWREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWREADY === 0 );
                    @( AWREADY );
                end
                while ( AWREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWREADY === 1 );
                    @( AWREADY );
                end
                while ( AWREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWUSER
    //     Wait for the specified change on wire <axi::AWUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWUSER === 0 );
                    @( AWUSER );
                end
                while ( AWUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWUSER === 1 );
                    @( AWUSER );
                end
                while ( AWUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWUSER_index1
    //     Wait for the specified change on wire <axi::AWUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWUSER[_this_dot_1] === 0 );
                    @( AWUSER[_this_dot_1] );
                end
                while ( AWUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWUSER[_this_dot_1] === 1 );
                    @( AWUSER[_this_dot_1] );
                end
                while ( AWUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARVALID
    //     Wait for the specified change on wire <axi::ARVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARVALID === 0 );
                    @( ARVALID );
                end
                while ( ARVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARVALID === 1 );
                    @( ARVALID );
                end
                while ( ARVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARADDR
    //     Wait for the specified change on wire <axi::ARADDR>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARADDR( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARADDR);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARADDR);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARADDR);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARADDR === 0 );
                    @( ARADDR );
                end
                while ( ARADDR !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARADDR === 1 );
                    @( ARADDR );
                end
                while ( ARADDR !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARADDR_index1
    //     Wait for the specified change on wire <axi::ARADDR>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARADDR_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARADDR[_this_dot_1] === 0 );
                    @( ARADDR[_this_dot_1] );
                end
                while ( ARADDR[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARADDR[_this_dot_1] === 1 );
                    @( ARADDR[_this_dot_1] );
                end
                while ( ARADDR[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLEN
    //     Wait for the specified change on wire <axi::ARLEN>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLEN( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLEN);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLEN);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLEN);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLEN === 0 );
                    @( ARLEN );
                end
                while ( ARLEN !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLEN === 1 );
                    @( ARLEN );
                end
                while ( ARLEN !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLEN_index1
    //     Wait for the specified change on wire <axi::ARLEN>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLEN_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLEN[_this_dot_1] === 0 );
                    @( ARLEN[_this_dot_1] );
                end
                while ( ARLEN[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLEN[_this_dot_1] === 1 );
                    @( ARLEN[_this_dot_1] );
                end
                while ( ARLEN[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARSIZE
    //     Wait for the specified change on wire <axi::ARSIZE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARSIZE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARSIZE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARSIZE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARSIZE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARSIZE === 0 );
                    @( ARSIZE );
                end
                while ( ARSIZE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARSIZE === 1 );
                    @( ARSIZE );
                end
                while ( ARSIZE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARSIZE_index1
    //     Wait for the specified change on wire <axi::ARSIZE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARSIZE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARSIZE[_this_dot_1] === 0 );
                    @( ARSIZE[_this_dot_1] );
                end
                while ( ARSIZE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARSIZE[_this_dot_1] === 1 );
                    @( ARSIZE[_this_dot_1] );
                end
                while ( ARSIZE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARBURST
    //     Wait for the specified change on wire <axi::ARBURST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARBURST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARBURST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARBURST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARBURST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARBURST === 0 );
                    @( ARBURST );
                end
                while ( ARBURST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARBURST === 1 );
                    @( ARBURST );
                end
                while ( ARBURST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARBURST_index1
    //     Wait for the specified change on wire <axi::ARBURST>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARBURST_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARBURST[_this_dot_1] === 0 );
                    @( ARBURST[_this_dot_1] );
                end
                while ( ARBURST[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARBURST[_this_dot_1] === 1 );
                    @( ARBURST[_this_dot_1] );
                end
                while ( ARBURST[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLOCK
    //     Wait for the specified change on wire <axi::ARLOCK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLOCK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLOCK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLOCK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLOCK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLOCK === 0 );
                    @( ARLOCK );
                end
                while ( ARLOCK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLOCK === 1 );
                    @( ARLOCK );
                end
                while ( ARLOCK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLOCK_index1
    //     Wait for the specified change on wire <axi::ARLOCK>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLOCK_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLOCK[_this_dot_1] === 0 );
                    @( ARLOCK[_this_dot_1] );
                end
                while ( ARLOCK[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLOCK[_this_dot_1] === 1 );
                    @( ARLOCK[_this_dot_1] );
                end
                while ( ARLOCK[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARCACHE
    //     Wait for the specified change on wire <axi::ARCACHE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARCACHE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARCACHE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARCACHE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARCACHE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARCACHE === 0 );
                    @( ARCACHE );
                end
                while ( ARCACHE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARCACHE === 1 );
                    @( ARCACHE );
                end
                while ( ARCACHE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARCACHE_index1
    //     Wait for the specified change on wire <axi::ARCACHE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARCACHE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARCACHE[_this_dot_1] === 0 );
                    @( ARCACHE[_this_dot_1] );
                end
                while ( ARCACHE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARCACHE[_this_dot_1] === 1 );
                    @( ARCACHE[_this_dot_1] );
                end
                while ( ARCACHE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARPROT
    //     Wait for the specified change on wire <axi::ARPROT>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARPROT( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARPROT);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARPROT);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARPROT);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARPROT === 0 );
                    @( ARPROT );
                end
                while ( ARPROT !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARPROT === 1 );
                    @( ARPROT );
                end
                while ( ARPROT !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARPROT_index1
    //     Wait for the specified change on wire <axi::ARPROT>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARPROT_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARPROT[_this_dot_1] === 0 );
                    @( ARPROT[_this_dot_1] );
                end
                while ( ARPROT[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARPROT[_this_dot_1] === 1 );
                    @( ARPROT[_this_dot_1] );
                end
                while ( ARPROT[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARID
    //     Wait for the specified change on wire <axi::ARID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARID === 0 );
                    @( ARID );
                end
                while ( ARID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARID === 1 );
                    @( ARID );
                end
                while ( ARID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARID_index1
    //     Wait for the specified change on wire <axi::ARID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARID[_this_dot_1] === 0 );
                    @( ARID[_this_dot_1] );
                end
                while ( ARID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARID[_this_dot_1] === 1 );
                    @( ARID[_this_dot_1] );
                end
                while ( ARID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARREADY
    //     Wait for the specified change on wire <axi::ARREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARREADY === 0 );
                    @( ARREADY );
                end
                while ( ARREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARREADY === 1 );
                    @( ARREADY );
                end
                while ( ARREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARUSER
    //     Wait for the specified change on wire <axi::ARUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARUSER === 0 );
                    @( ARUSER );
                end
                while ( ARUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARUSER === 1 );
                    @( ARUSER );
                end
                while ( ARUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARUSER_index1
    //     Wait for the specified change on wire <axi::ARUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARUSER[_this_dot_1] === 0 );
                    @( ARUSER[_this_dot_1] );
                end
                while ( ARUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARUSER[_this_dot_1] === 1 );
                    @( ARUSER[_this_dot_1] );
                end
                while ( ARUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RVALID
    //     Wait for the specified change on wire <axi::RVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RVALID === 0 );
                    @( RVALID );
                end
                while ( RVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RVALID === 1 );
                    @( RVALID );
                end
                while ( RVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RLAST
    //     Wait for the specified change on wire <axi::RLAST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RLAST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RLAST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RLAST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RLAST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RLAST === 0 );
                    @( RLAST );
                end
                while ( RLAST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RLAST === 1 );
                    @( RLAST );
                end
                while ( RLAST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RDATA
    //     Wait for the specified change on wire <axi::RDATA>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RDATA( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RDATA);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RDATA);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RDATA);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RDATA === 0 );
                    @( RDATA );
                end
                while ( RDATA !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RDATA === 1 );
                    @( RDATA );
                end
                while ( RDATA !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RDATA_index1
    //     Wait for the specified change on wire <axi::RDATA>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RDATA_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RDATA[_this_dot_1] === 0 );
                    @( RDATA[_this_dot_1] );
                end
                while ( RDATA[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RDATA[_this_dot_1] === 1 );
                    @( RDATA[_this_dot_1] );
                end
                while ( RDATA[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RRESP
    //     Wait for the specified change on wire <axi::RRESP>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RRESP( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RRESP);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RRESP);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RRESP);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RRESP === 0 );
                    @( RRESP );
                end
                while ( RRESP !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RRESP === 1 );
                    @( RRESP );
                end
                while ( RRESP !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RRESP_index1
    //     Wait for the specified change on wire <axi::RRESP>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RRESP_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RRESP[_this_dot_1] === 0 );
                    @( RRESP[_this_dot_1] );
                end
                while ( RRESP[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RRESP[_this_dot_1] === 1 );
                    @( RRESP[_this_dot_1] );
                end
                while ( RRESP[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RID
    //     Wait for the specified change on wire <axi::RID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RID === 0 );
                    @( RID );
                end
                while ( RID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RID === 1 );
                    @( RID );
                end
                while ( RID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RID_index1
    //     Wait for the specified change on wire <axi::RID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RID[_this_dot_1] === 0 );
                    @( RID[_this_dot_1] );
                end
                while ( RID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RID[_this_dot_1] === 1 );
                    @( RID[_this_dot_1] );
                end
                while ( RID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RREADY
    //     Wait for the specified change on wire <axi::RREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RREADY === 0 );
                    @( RREADY );
                end
                while ( RREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RREADY === 1 );
                    @( RREADY );
                end
                while ( RREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RUSER
    //     Wait for the specified change on wire <axi::RUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RUSER === 0 );
                    @( RUSER );
                end
                while ( RUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RUSER === 1 );
                    @( RUSER );
                end
                while ( RUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RUSER_index1
    //     Wait for the specified change on wire <axi::RUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RUSER[_this_dot_1] === 0 );
                    @( RUSER[_this_dot_1] );
                end
                while ( RUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RUSER[_this_dot_1] === 1 );
                    @( RUSER[_this_dot_1] );
                end
                while ( RUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WVALID
    //     Wait for the specified change on wire <axi::WVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WVALID === 0 );
                    @( WVALID );
                end
                while ( WVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WVALID === 1 );
                    @( WVALID );
                end
                while ( WVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WLAST
    //     Wait for the specified change on wire <axi::WLAST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WLAST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WLAST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WLAST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WLAST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WLAST === 0 );
                    @( WLAST );
                end
                while ( WLAST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WLAST === 1 );
                    @( WLAST );
                end
                while ( WLAST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WDATA
    //     Wait for the specified change on wire <axi::WDATA>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WDATA( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WDATA);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WDATA);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WDATA);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WDATA === 0 );
                    @( WDATA );
                end
                while ( WDATA !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WDATA === 1 );
                    @( WDATA );
                end
                while ( WDATA !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WDATA_index1
    //     Wait for the specified change on wire <axi::WDATA>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WDATA_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WDATA[_this_dot_1] === 0 );
                    @( WDATA[_this_dot_1] );
                end
                while ( WDATA[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WDATA[_this_dot_1] === 1 );
                    @( WDATA[_this_dot_1] );
                end
                while ( WDATA[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WSTRB
    //     Wait for the specified change on wire <axi::WSTRB>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WSTRB( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WSTRB);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WSTRB);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WSTRB);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WSTRB === 0 );
                    @( WSTRB );
                end
                while ( WSTRB !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WSTRB === 1 );
                    @( WSTRB );
                end
                while ( WSTRB !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WSTRB_index1
    //     Wait for the specified change on wire <axi::WSTRB>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WSTRB_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WSTRB[_this_dot_1] === 0 );
                    @( WSTRB[_this_dot_1] );
                end
                while ( WSTRB[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WSTRB[_this_dot_1] === 1 );
                    @( WSTRB[_this_dot_1] );
                end
                while ( WSTRB[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WID
    //     Wait for the specified change on wire <axi::WID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WID === 0 );
                    @( WID );
                end
                while ( WID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WID === 1 );
                    @( WID );
                end
                while ( WID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WID_index1
    //     Wait for the specified change on wire <axi::WID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WID[_this_dot_1] === 0 );
                    @( WID[_this_dot_1] );
                end
                while ( WID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WID[_this_dot_1] === 1 );
                    @( WID[_this_dot_1] );
                end
                while ( WID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WREADY
    //     Wait for the specified change on wire <axi::WREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WREADY === 0 );
                    @( WREADY );
                end
                while ( WREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WREADY === 1 );
                    @( WREADY );
                end
                while ( WREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WUSER
    //     Wait for the specified change on wire <axi::WUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WUSER === 0 );
                    @( WUSER );
                end
                while ( WUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WUSER === 1 );
                    @( WUSER );
                end
                while ( WUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WUSER_index1
    //     Wait for the specified change on wire <axi::WUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WUSER[_this_dot_1] === 0 );
                    @( WUSER[_this_dot_1] );
                end
                while ( WUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WUSER[_this_dot_1] === 1 );
                    @( WUSER[_this_dot_1] );
                end
                while ( WUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BVALID
    //     Wait for the specified change on wire <axi::BVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BVALID === 0 );
                    @( BVALID );
                end
                while ( BVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BVALID === 1 );
                    @( BVALID );
                end
                while ( BVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BRESP
    //     Wait for the specified change on wire <axi::BRESP>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BRESP( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BRESP);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BRESP);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BRESP);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BRESP === 0 );
                    @( BRESP );
                end
                while ( BRESP !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BRESP === 1 );
                    @( BRESP );
                end
                while ( BRESP !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BRESP_index1
    //     Wait for the specified change on wire <axi::BRESP>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BRESP_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BRESP[_this_dot_1] === 0 );
                    @( BRESP[_this_dot_1] );
                end
                while ( BRESP[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BRESP[_this_dot_1] === 1 );
                    @( BRESP[_this_dot_1] );
                end
                while ( BRESP[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BID
    //     Wait for the specified change on wire <axi::BID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BID === 0 );
                    @( BID );
                end
                while ( BID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BID === 1 );
                    @( BID );
                end
                while ( BID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BID_index1
    //     Wait for the specified change on wire <axi::BID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BID[_this_dot_1] === 0 );
                    @( BID[_this_dot_1] );
                end
                while ( BID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BID[_this_dot_1] === 1 );
                    @( BID[_this_dot_1] );
                end
                while ( BID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BREADY
    //     Wait for the specified change on wire <axi::BREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BREADY === 0 );
                    @( BREADY );
                end
                while ( BREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BREADY === 1 );
                    @( BREADY );
                end
                while ( BREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BUSER
    //     Wait for the specified change on wire <axi::BUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BUSER === 0 );
                    @( BUSER );
                end
                while ( BUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BUSER === 1 );
                    @( BUSER );
                end
                while ( BUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BUSER_index1
    //     Wait for the specified change on wire <axi::BUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BUSER[_this_dot_1] === 0 );
                    @( BUSER[_this_dot_1] );
                end
                while ( BUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BUSER[_this_dot_1] === 1 );
                    @( BUSER[_this_dot_1] );
                end
                while ( BUSER[_this_dot_1] !== 0 );
            end
        end
    endtask

    //-------------------------------------------------------------------------
    // Tasks/functions to set/get wires
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- set_ACLK
    //-------------------------------------------------------------------------
    //     Set the value of wire <ACLK>.
    //
    // Parameters:
    //     ACLK_param - The value to set onto wire <ACLK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ACLK( logic ACLK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ACLK = ACLK_param;
        else
            m_ACLK <= ACLK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ACLK
    //-------------------------------------------------------------------------
    //     Get the value of wire <ACLK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ACLK>.
    //
    function automatic logic get_ACLK(  );
        return ACLK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARESETn
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARESETn>.
    //
    // Parameters:
    //     ARESETn_param - The value to set onto wire <ARESETn>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARESETn( logic ARESETn_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARESETn = ARESETn_param;
        else
            m_ARESETn <= ARESETn_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARESETn
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARESETn>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARESETn>.
    //
    function automatic logic get_ARESETn(  );
        return ARESETn;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWVALID>.
    //
    // Parameters:
    //     AWVALID_param - The value to set onto wire <AWVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWVALID( logic AWVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWVALID = AWVALID_param;
        else
            m_AWVALID <= AWVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWVALID>.
    //
    function automatic logic get_AWVALID(  );
        return AWVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWADDR
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWADDR>.
    //
    // Parameters:
    //     AWADDR_param - The value to set onto wire <AWADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWADDR( logic [((AXI_ADDRESS_WIDTH) - 1):0]  AWADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWADDR = AWADDR_param;
        else
            m_AWADDR <= AWADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWADDR_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWADDR_param - The value to set onto wire <AWADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWADDR_index1( int _this_dot_1, logic  AWADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWADDR[_this_dot_1] = AWADDR_param;
        else
            m_AWADDR[_this_dot_1] <= AWADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWADDR
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWADDR>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWADDR>.
    //
    function automatic logic [((AXI_ADDRESS_WIDTH) - 1):0]   get_AWADDR(  );
        return AWADDR;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWADDR_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWADDR>.
    //
    function automatic logic   get_AWADDR_index1( int _this_dot_1 );
        return AWADDR[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWLEN
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWLEN>.
    //
    // Parameters:
    //     AWLEN_param - The value to set onto wire <AWLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLEN( logic [3:0] AWLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLEN = AWLEN_param;
        else
            m_AWLEN <= AWLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWLEN_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWLEN_param - The value to set onto wire <AWLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLEN_index1( int _this_dot_1, logic  AWLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLEN[_this_dot_1] = AWLEN_param;
        else
            m_AWLEN[_this_dot_1] <= AWLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWLEN
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWLEN>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWLEN>.
    //
    function automatic logic [3:0]  get_AWLEN(  );
        return AWLEN;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWLEN_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWLEN>.
    //
    function automatic logic   get_AWLEN_index1( int _this_dot_1 );
        return AWLEN[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWSIZE
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWSIZE>.
    //
    // Parameters:
    //     AWSIZE_param - The value to set onto wire <AWSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWSIZE( logic [2:0] AWSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWSIZE = AWSIZE_param;
        else
            m_AWSIZE <= AWSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWSIZE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWSIZE_param - The value to set onto wire <AWSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWSIZE_index1( int _this_dot_1, logic  AWSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWSIZE[_this_dot_1] = AWSIZE_param;
        else
            m_AWSIZE[_this_dot_1] <= AWSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWSIZE
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWSIZE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWSIZE>.
    //
    function automatic logic [2:0]  get_AWSIZE(  );
        return AWSIZE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWSIZE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWSIZE>.
    //
    function automatic logic   get_AWSIZE_index1( int _this_dot_1 );
        return AWSIZE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWBURST
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWBURST>.
    //
    // Parameters:
    //     AWBURST_param - The value to set onto wire <AWBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWBURST( logic [1:0] AWBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWBURST = AWBURST_param;
        else
            m_AWBURST <= AWBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWBURST_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWBURST_param - The value to set onto wire <AWBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWBURST_index1( int _this_dot_1, logic  AWBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWBURST[_this_dot_1] = AWBURST_param;
        else
            m_AWBURST[_this_dot_1] <= AWBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWBURST
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWBURST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWBURST>.
    //
    function automatic logic [1:0]  get_AWBURST(  );
        return AWBURST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWBURST_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWBURST>.
    //
    function automatic logic   get_AWBURST_index1( int _this_dot_1 );
        return AWBURST[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWLOCK
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWLOCK>.
    //
    // Parameters:
    //     AWLOCK_param - The value to set onto wire <AWLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLOCK( logic [1:0] AWLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLOCK = AWLOCK_param;
        else
            m_AWLOCK <= AWLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWLOCK_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWLOCK_param - The value to set onto wire <AWLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLOCK_index1( int _this_dot_1, logic  AWLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLOCK[_this_dot_1] = AWLOCK_param;
        else
            m_AWLOCK[_this_dot_1] <= AWLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWLOCK
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWLOCK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWLOCK>.
    //
    function automatic logic [1:0]  get_AWLOCK(  );
        return AWLOCK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWLOCK_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWLOCK>.
    //
    function automatic logic   get_AWLOCK_index1( int _this_dot_1 );
        return AWLOCK[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWCACHE
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWCACHE>.
    //
    // Parameters:
    //     AWCACHE_param - The value to set onto wire <AWCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWCACHE( logic [3:0] AWCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWCACHE = AWCACHE_param;
        else
            m_AWCACHE <= AWCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWCACHE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWCACHE_param - The value to set onto wire <AWCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWCACHE_index1( int _this_dot_1, logic  AWCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWCACHE[_this_dot_1] = AWCACHE_param;
        else
            m_AWCACHE[_this_dot_1] <= AWCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWCACHE
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWCACHE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWCACHE>.
    //
    function automatic logic [3:0]  get_AWCACHE(  );
        return AWCACHE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWCACHE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWCACHE>.
    //
    function automatic logic   get_AWCACHE_index1( int _this_dot_1 );
        return AWCACHE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWPROT
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWPROT>.
    //
    // Parameters:
    //     AWPROT_param - The value to set onto wire <AWPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWPROT( logic [2:0] AWPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWPROT = AWPROT_param;
        else
            m_AWPROT <= AWPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWPROT_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWPROT_param - The value to set onto wire <AWPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWPROT_index1( int _this_dot_1, logic  AWPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWPROT[_this_dot_1] = AWPROT_param;
        else
            m_AWPROT[_this_dot_1] <= AWPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWPROT
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWPROT>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWPROT>.
    //
    function automatic logic [2:0]  get_AWPROT(  );
        return AWPROT;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWPROT_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWPROT>.
    //
    function automatic logic   get_AWPROT_index1( int _this_dot_1 );
        return AWPROT[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWID
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWID>.
    //
    // Parameters:
    //     AWID_param - The value to set onto wire <AWID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWID( logic [((AXI_ID_WIDTH) - 1):0]  AWID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWID = AWID_param;
        else
            m_AWID <= AWID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWID_param - The value to set onto wire <AWID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWID_index1( int _this_dot_1, logic  AWID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWID[_this_dot_1] = AWID_param;
        else
            m_AWID[_this_dot_1] <= AWID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWID
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_AWID(  );
        return AWID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWID>.
    //
    function automatic logic   get_AWID_index1( int _this_dot_1 );
        return AWID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWREADY>.
    //
    // Parameters:
    //     AWREADY_param - The value to set onto wire <AWREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWREADY( logic AWREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWREADY = AWREADY_param;
        else
            m_AWREADY <= AWREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWREADY>.
    //
    function automatic logic get_AWREADY(  );
        return AWREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWUSER>.
    //
    // Parameters:
    //     AWUSER_param - The value to set onto wire <AWUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWUSER( logic [7:0] AWUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWUSER = AWUSER_param;
        else
            m_AWUSER <= AWUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWUSER_param - The value to set onto wire <AWUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWUSER_index1( int _this_dot_1, logic  AWUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWUSER[_this_dot_1] = AWUSER_param;
        else
            m_AWUSER[_this_dot_1] <= AWUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWUSER>.
    //
    function automatic logic [7:0]  get_AWUSER(  );
        return AWUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWUSER>.
    //
    function automatic logic   get_AWUSER_index1( int _this_dot_1 );
        return AWUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARVALID>.
    //
    // Parameters:
    //     ARVALID_param - The value to set onto wire <ARVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARVALID( logic ARVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARVALID = ARVALID_param;
        else
            m_ARVALID <= ARVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARVALID>.
    //
    function automatic logic get_ARVALID(  );
        return ARVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARADDR
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARADDR>.
    //
    // Parameters:
    //     ARADDR_param - The value to set onto wire <ARADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARADDR( logic [((AXI_ADDRESS_WIDTH) - 1):0]  ARADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARADDR = ARADDR_param;
        else
            m_ARADDR <= ARADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARADDR_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARADDR_param - The value to set onto wire <ARADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARADDR_index1( int _this_dot_1, logic  ARADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARADDR[_this_dot_1] = ARADDR_param;
        else
            m_ARADDR[_this_dot_1] <= ARADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARADDR
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARADDR>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARADDR>.
    //
    function automatic logic [((AXI_ADDRESS_WIDTH) - 1):0]   get_ARADDR(  );
        return ARADDR;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARADDR_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARADDR>.
    //
    function automatic logic   get_ARADDR_index1( int _this_dot_1 );
        return ARADDR[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARLEN
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARLEN>.
    //
    // Parameters:
    //     ARLEN_param - The value to set onto wire <ARLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLEN( logic [3:0] ARLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLEN = ARLEN_param;
        else
            m_ARLEN <= ARLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARLEN_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARLEN_param - The value to set onto wire <ARLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLEN_index1( int _this_dot_1, logic  ARLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLEN[_this_dot_1] = ARLEN_param;
        else
            m_ARLEN[_this_dot_1] <= ARLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARLEN
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARLEN>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARLEN>.
    //
    function automatic logic [3:0]  get_ARLEN(  );
        return ARLEN;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARLEN_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARLEN>.
    //
    function automatic logic   get_ARLEN_index1( int _this_dot_1 );
        return ARLEN[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARSIZE
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARSIZE>.
    //
    // Parameters:
    //     ARSIZE_param - The value to set onto wire <ARSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARSIZE( logic [2:0] ARSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARSIZE = ARSIZE_param;
        else
            m_ARSIZE <= ARSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARSIZE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARSIZE_param - The value to set onto wire <ARSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARSIZE_index1( int _this_dot_1, logic  ARSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARSIZE[_this_dot_1] = ARSIZE_param;
        else
            m_ARSIZE[_this_dot_1] <= ARSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARSIZE
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARSIZE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARSIZE>.
    //
    function automatic logic [2:0]  get_ARSIZE(  );
        return ARSIZE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARSIZE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARSIZE>.
    //
    function automatic logic   get_ARSIZE_index1( int _this_dot_1 );
        return ARSIZE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARBURST
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARBURST>.
    //
    // Parameters:
    //     ARBURST_param - The value to set onto wire <ARBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARBURST( logic [1:0] ARBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARBURST = ARBURST_param;
        else
            m_ARBURST <= ARBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARBURST_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARBURST_param - The value to set onto wire <ARBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARBURST_index1( int _this_dot_1, logic  ARBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARBURST[_this_dot_1] = ARBURST_param;
        else
            m_ARBURST[_this_dot_1] <= ARBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARBURST
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARBURST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARBURST>.
    //
    function automatic logic [1:0]  get_ARBURST(  );
        return ARBURST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARBURST_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARBURST>.
    //
    function automatic logic   get_ARBURST_index1( int _this_dot_1 );
        return ARBURST[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARLOCK
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARLOCK>.
    //
    // Parameters:
    //     ARLOCK_param - The value to set onto wire <ARLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLOCK( logic [1:0] ARLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLOCK = ARLOCK_param;
        else
            m_ARLOCK <= ARLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARLOCK_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARLOCK_param - The value to set onto wire <ARLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLOCK_index1( int _this_dot_1, logic  ARLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLOCK[_this_dot_1] = ARLOCK_param;
        else
            m_ARLOCK[_this_dot_1] <= ARLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARLOCK
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARLOCK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARLOCK>.
    //
    function automatic logic [1:0]  get_ARLOCK(  );
        return ARLOCK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARLOCK_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARLOCK>.
    //
    function automatic logic   get_ARLOCK_index1( int _this_dot_1 );
        return ARLOCK[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARCACHE
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARCACHE>.
    //
    // Parameters:
    //     ARCACHE_param - The value to set onto wire <ARCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARCACHE( logic [3:0] ARCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARCACHE = ARCACHE_param;
        else
            m_ARCACHE <= ARCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARCACHE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARCACHE_param - The value to set onto wire <ARCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARCACHE_index1( int _this_dot_1, logic  ARCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARCACHE[_this_dot_1] = ARCACHE_param;
        else
            m_ARCACHE[_this_dot_1] <= ARCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARCACHE
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARCACHE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARCACHE>.
    //
    function automatic logic [3:0]  get_ARCACHE(  );
        return ARCACHE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARCACHE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARCACHE>.
    //
    function automatic logic   get_ARCACHE_index1( int _this_dot_1 );
        return ARCACHE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARPROT
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARPROT>.
    //
    // Parameters:
    //     ARPROT_param - The value to set onto wire <ARPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARPROT( logic [2:0] ARPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARPROT = ARPROT_param;
        else
            m_ARPROT <= ARPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARPROT_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARPROT_param - The value to set onto wire <ARPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARPROT_index1( int _this_dot_1, logic  ARPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARPROT[_this_dot_1] = ARPROT_param;
        else
            m_ARPROT[_this_dot_1] <= ARPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARPROT
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARPROT>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARPROT>.
    //
    function automatic logic [2:0]  get_ARPROT(  );
        return ARPROT;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARPROT_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARPROT>.
    //
    function automatic logic   get_ARPROT_index1( int _this_dot_1 );
        return ARPROT[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARID
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARID>.
    //
    // Parameters:
    //     ARID_param - The value to set onto wire <ARID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARID( logic [((AXI_ID_WIDTH) - 1):0]  ARID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARID = ARID_param;
        else
            m_ARID <= ARID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARID_param - The value to set onto wire <ARID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARID_index1( int _this_dot_1, logic  ARID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARID[_this_dot_1] = ARID_param;
        else
            m_ARID[_this_dot_1] <= ARID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARID
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_ARID(  );
        return ARID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARID>.
    //
    function automatic logic   get_ARID_index1( int _this_dot_1 );
        return ARID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARREADY>.
    //
    // Parameters:
    //     ARREADY_param - The value to set onto wire <ARREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARREADY( logic ARREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARREADY = ARREADY_param;
        else
            m_ARREADY <= ARREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARREADY>.
    //
    function automatic logic get_ARREADY(  );
        return ARREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARUSER>.
    //
    // Parameters:
    //     ARUSER_param - The value to set onto wire <ARUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARUSER( logic [7:0] ARUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARUSER = ARUSER_param;
        else
            m_ARUSER <= ARUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARUSER_param - The value to set onto wire <ARUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARUSER_index1( int _this_dot_1, logic  ARUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARUSER[_this_dot_1] = ARUSER_param;
        else
            m_ARUSER[_this_dot_1] <= ARUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARUSER>.
    //
    function automatic logic [7:0]  get_ARUSER(  );
        return ARUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARUSER>.
    //
    function automatic logic   get_ARUSER_index1( int _this_dot_1 );
        return ARUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <RVALID>.
    //
    // Parameters:
    //     RVALID_param - The value to set onto wire <RVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RVALID( logic RVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RVALID = RVALID_param;
        else
            m_RVALID <= RVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <RVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RVALID>.
    //
    function automatic logic get_RVALID(  );
        return RVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RLAST
    //-------------------------------------------------------------------------
    //     Set the value of wire <RLAST>.
    //
    // Parameters:
    //     RLAST_param - The value to set onto wire <RLAST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RLAST( logic RLAST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RLAST = RLAST_param;
        else
            m_RLAST <= RLAST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RLAST
    //-------------------------------------------------------------------------
    //     Get the value of wire <RLAST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RLAST>.
    //
    function automatic logic get_RLAST(  );
        return RLAST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RDATA
    //-------------------------------------------------------------------------
    //     Set the value of wire <RDATA>.
    //
    // Parameters:
    //     RDATA_param - The value to set onto wire <RDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RDATA( logic [((AXI_RDATA_WIDTH) - 1):0]  RDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RDATA = RDATA_param;
        else
            m_RDATA <= RDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RDATA_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RDATA_param - The value to set onto wire <RDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RDATA_index1( int _this_dot_1, logic  RDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RDATA[_this_dot_1] = RDATA_param;
        else
            m_RDATA[_this_dot_1] <= RDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RDATA
    //-------------------------------------------------------------------------
    //     Get the value of wire <RDATA>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RDATA>.
    //
    function automatic logic [((AXI_RDATA_WIDTH) - 1):0]   get_RDATA(  );
        return RDATA;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RDATA_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RDATA>.
    //
    function automatic logic   get_RDATA_index1( int _this_dot_1 );
        return RDATA[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RRESP
    //-------------------------------------------------------------------------
    //     Set the value of wire <RRESP>.
    //
    // Parameters:
    //     RRESP_param - The value to set onto wire <RRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RRESP( logic [1:0] RRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RRESP = RRESP_param;
        else
            m_RRESP <= RRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RRESP_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RRESP_param - The value to set onto wire <RRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RRESP_index1( int _this_dot_1, logic  RRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RRESP[_this_dot_1] = RRESP_param;
        else
            m_RRESP[_this_dot_1] <= RRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RRESP
    //-------------------------------------------------------------------------
    //     Get the value of wire <RRESP>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RRESP>.
    //
    function automatic logic [1:0]  get_RRESP(  );
        return RRESP;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RRESP_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RRESP>.
    //
    function automatic logic   get_RRESP_index1( int _this_dot_1 );
        return RRESP[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RID
    //-------------------------------------------------------------------------
    //     Set the value of wire <RID>.
    //
    // Parameters:
    //     RID_param - The value to set onto wire <RID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RID( logic [((AXI_ID_WIDTH) - 1):0]  RID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RID = RID_param;
        else
            m_RID <= RID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RID_param - The value to set onto wire <RID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RID_index1( int _this_dot_1, logic  RID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RID[_this_dot_1] = RID_param;
        else
            m_RID[_this_dot_1] <= RID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RID
    //-------------------------------------------------------------------------
    //     Get the value of wire <RID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_RID(  );
        return RID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RID>.
    //
    function automatic logic   get_RID_index1( int _this_dot_1 );
        return RID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <RREADY>.
    //
    // Parameters:
    //     RREADY_param - The value to set onto wire <RREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RREADY( logic RREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RREADY = RREADY_param;
        else
            m_RREADY <= RREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <RREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RREADY>.
    //
    function automatic logic get_RREADY(  );
        return RREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <RUSER>.
    //
    // Parameters:
    //     RUSER_param - The value to set onto wire <RUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RUSER( logic [7:0] RUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RUSER = RUSER_param;
        else
            m_RUSER <= RUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RUSER_param - The value to set onto wire <RUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RUSER_index1( int _this_dot_1, logic  RUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RUSER[_this_dot_1] = RUSER_param;
        else
            m_RUSER[_this_dot_1] <= RUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <RUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RUSER>.
    //
    function automatic logic [7:0]  get_RUSER(  );
        return RUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RUSER>.
    //
    function automatic logic   get_RUSER_index1( int _this_dot_1 );
        return RUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <WVALID>.
    //
    // Parameters:
    //     WVALID_param - The value to set onto wire <WVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WVALID( logic WVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WVALID = WVALID_param;
        else
            m_WVALID <= WVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <WVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WVALID>.
    //
    function automatic logic get_WVALID(  );
        return WVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WLAST
    //-------------------------------------------------------------------------
    //     Set the value of wire <WLAST>.
    //
    // Parameters:
    //     WLAST_param - The value to set onto wire <WLAST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WLAST( logic WLAST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WLAST = WLAST_param;
        else
            m_WLAST <= WLAST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WLAST
    //-------------------------------------------------------------------------
    //     Get the value of wire <WLAST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WLAST>.
    //
    function automatic logic get_WLAST(  );
        return WLAST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WDATA
    //-------------------------------------------------------------------------
    //     Set the value of wire <WDATA>.
    //
    // Parameters:
    //     WDATA_param - The value to set onto wire <WDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WDATA( logic [((AXI_WDATA_WIDTH) - 1):0]  WDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WDATA = WDATA_param;
        else
            m_WDATA <= WDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WDATA_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WDATA_param - The value to set onto wire <WDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WDATA_index1( int _this_dot_1, logic  WDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WDATA[_this_dot_1] = WDATA_param;
        else
            m_WDATA[_this_dot_1] <= WDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WDATA
    //-------------------------------------------------------------------------
    //     Get the value of wire <WDATA>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WDATA>.
    //
    function automatic logic [((AXI_WDATA_WIDTH) - 1):0]   get_WDATA(  );
        return WDATA;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WDATA_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WDATA>.
    //
    function automatic logic   get_WDATA_index1( int _this_dot_1 );
        return WDATA[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WSTRB
    //-------------------------------------------------------------------------
    //     Set the value of wire <WSTRB>.
    //
    // Parameters:
    //     WSTRB_param - The value to set onto wire <WSTRB>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WSTRB( logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  WSTRB_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WSTRB = WSTRB_param;
        else
            m_WSTRB <= WSTRB_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WSTRB_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WSTRB>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WSTRB_param - The value to set onto wire <WSTRB>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WSTRB_index1( int _this_dot_1, logic  WSTRB_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WSTRB[_this_dot_1] = WSTRB_param;
        else
            m_WSTRB[_this_dot_1] <= WSTRB_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WSTRB
    //-------------------------------------------------------------------------
    //     Get the value of wire <WSTRB>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WSTRB>.
    //
    function automatic logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]   get_WSTRB(  );
        return WSTRB;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WSTRB_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WSTRB>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WSTRB>.
    //
    function automatic logic   get_WSTRB_index1( int _this_dot_1 );
        return WSTRB[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WID
    //-------------------------------------------------------------------------
    //     Set the value of wire <WID>.
    //
    // Parameters:
    //     WID_param - The value to set onto wire <WID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WID( logic [((AXI_ID_WIDTH) - 1):0]  WID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WID = WID_param;
        else
            m_WID <= WID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WID_param - The value to set onto wire <WID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WID_index1( int _this_dot_1, logic  WID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WID[_this_dot_1] = WID_param;
        else
            m_WID[_this_dot_1] <= WID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WID
    //-------------------------------------------------------------------------
    //     Get the value of wire <WID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_WID(  );
        return WID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WID>.
    //
    function automatic logic   get_WID_index1( int _this_dot_1 );
        return WID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <WREADY>.
    //
    // Parameters:
    //     WREADY_param - The value to set onto wire <WREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WREADY( logic WREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WREADY = WREADY_param;
        else
            m_WREADY <= WREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <WREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WREADY>.
    //
    function automatic logic get_WREADY(  );
        return WREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <WUSER>.
    //
    // Parameters:
    //     WUSER_param - The value to set onto wire <WUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WUSER( logic [7:0] WUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WUSER = WUSER_param;
        else
            m_WUSER <= WUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WUSER_param - The value to set onto wire <WUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WUSER_index1( int _this_dot_1, logic  WUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WUSER[_this_dot_1] = WUSER_param;
        else
            m_WUSER[_this_dot_1] <= WUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <WUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WUSER>.
    //
    function automatic logic [7:0]  get_WUSER(  );
        return WUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WUSER>.
    //
    function automatic logic   get_WUSER_index1( int _this_dot_1 );
        return WUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <BVALID>.
    //
    // Parameters:
    //     BVALID_param - The value to set onto wire <BVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BVALID( logic BVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BVALID = BVALID_param;
        else
            m_BVALID <= BVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <BVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BVALID>.
    //
    function automatic logic get_BVALID(  );
        return BVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BRESP
    //-------------------------------------------------------------------------
    //     Set the value of wire <BRESP>.
    //
    // Parameters:
    //     BRESP_param - The value to set onto wire <BRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BRESP( logic [1:0] BRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BRESP = BRESP_param;
        else
            m_BRESP <= BRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BRESP_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BRESP_param - The value to set onto wire <BRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BRESP_index1( int _this_dot_1, logic  BRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BRESP[_this_dot_1] = BRESP_param;
        else
            m_BRESP[_this_dot_1] <= BRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BRESP
    //-------------------------------------------------------------------------
    //     Get the value of wire <BRESP>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BRESP>.
    //
    function automatic logic [1:0]  get_BRESP(  );
        return BRESP;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BRESP_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BRESP>.
    //
    function automatic logic   get_BRESP_index1( int _this_dot_1 );
        return BRESP[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BID
    //-------------------------------------------------------------------------
    //     Set the value of wire <BID>.
    //
    // Parameters:
    //     BID_param - The value to set onto wire <BID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BID( logic [((AXI_ID_WIDTH) - 1):0]  BID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BID = BID_param;
        else
            m_BID <= BID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BID_param - The value to set onto wire <BID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BID_index1( int _this_dot_1, logic  BID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BID[_this_dot_1] = BID_param;
        else
            m_BID[_this_dot_1] <= BID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BID
    //-------------------------------------------------------------------------
    //     Get the value of wire <BID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_BID(  );
        return BID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BID>.
    //
    function automatic logic   get_BID_index1( int _this_dot_1 );
        return BID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <BREADY>.
    //
    // Parameters:
    //     BREADY_param - The value to set onto wire <BREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BREADY( logic BREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BREADY = BREADY_param;
        else
            m_BREADY <= BREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <BREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BREADY>.
    //
    function automatic logic get_BREADY(  );
        return BREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <BUSER>.
    //
    // Parameters:
    //     BUSER_param - The value to set onto wire <BUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BUSER( logic [7:0] BUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BUSER = BUSER_param;
        else
            m_BUSER <= BUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BUSER_param - The value to set onto wire <BUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BUSER_index1( int _this_dot_1, logic  BUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BUSER[_this_dot_1] = BUSER_param;
        else
            m_BUSER[_this_dot_1] <= BUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <BUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BUSER>.
    //
    function automatic logic [7:0]  get_BUSER(  );
        return BUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BUSER>.
    //
    function automatic logic   get_BUSER_index1( int _this_dot_1 );
        return BUSER[_this_dot_1];
    endfunction

    //-------------------------------------------------------------------------
    // Tasks to wait for a change to a global variable with read access
    //-------------------------------------------------------------------------


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_write_ctrl_to_data_mintime
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_write_ctrl_to_data_mintime>.
    //
    task automatic wait_for_config_write_ctrl_to_data_mintime(  );
        begin
            @( config_write_ctrl_to_data_mintime );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_master_write_delay
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_master_write_delay>.
    //
    task automatic wait_for_config_master_write_delay(  );
        begin
            @( config_master_write_delay );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_all_assertions
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_all_assertions>.
    //
    task automatic wait_for_config_enable_all_assertions(  );
        begin
            @( config_enable_all_assertions );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_assertion
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_assertion>.
    //
    task automatic wait_for_config_enable_assertion(  );
        begin
            @( config_enable_assertion );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_assertion_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_enable_assertion_index1( input int _this_dot_1 );
        begin
            @( config_enable_assertion[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_start_addr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_start_addr>.
    //
    task automatic wait_for_config_slave_start_addr(  );
        begin
            @( config_slave_start_addr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_start_addr_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_slave_start_addr_index1( input int _this_dot_1 );
        begin
            @( config_slave_start_addr[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_end_addr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_end_addr>.
    //
    task automatic wait_for_config_slave_end_addr(  );
        begin
            @( config_slave_end_addr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_end_addr_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_slave_end_addr_index1( input int _this_dot_1 );
        begin
            @( config_slave_end_addr[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_support_exclusive_access
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_support_exclusive_access>.
    //
    task automatic wait_for_config_support_exclusive_access(  );
        begin
            @( config_support_exclusive_access );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_read_data_reordering_depth
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_read_data_reordering_depth>.
    //
    task automatic wait_for_config_read_data_reordering_depth(  );
        begin
            @( config_read_data_reordering_depth );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_transaction_time_factor
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_transaction_time_factor>.
    //
    task automatic wait_for_config_max_transaction_time_factor(  );
        begin
            @( config_max_transaction_time_factor );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_timeout_max_data_transfer
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_timeout_max_data_transfer>.
    //
    task automatic wait_for_config_timeout_max_data_transfer(  );
        begin
            @( config_timeout_max_data_transfer );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_burst_timeout_factor
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_burst_timeout_factor>.
    //
    task automatic wait_for_config_burst_timeout_factor(  );
        begin
            @( config_burst_timeout_factor );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_AWVALID_assertion_to_AWREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    task automatic wait_for_config_max_latency_AWVALID_assertion_to_AWREADY(  );
        begin
            @( config_max_latency_AWVALID_assertion_to_AWREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_ARVALID_assertion_to_ARREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    task automatic wait_for_config_max_latency_ARVALID_assertion_to_ARREADY(  );
        begin
            @( config_max_latency_ARVALID_assertion_to_ARREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_RVALID_assertion_to_RREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_RVALID_assertion_to_RREADY>.
    //
    task automatic wait_for_config_max_latency_RVALID_assertion_to_RREADY(  );
        begin
            @( config_max_latency_RVALID_assertion_to_RREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_BVALID_assertion_to_BREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_BVALID_assertion_to_BREADY>.
    //
    task automatic wait_for_config_max_latency_BVALID_assertion_to_BREADY(  );
        begin
            @( config_max_latency_BVALID_assertion_to_BREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_WVALID_assertion_to_WREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_WVALID_assertion_to_WREADY>.
    //
    task automatic wait_for_config_max_latency_WVALID_assertion_to_WREADY(  );
        begin
            @( config_max_latency_WVALID_assertion_to_WREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_master_error_position
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_master_error_position>.
    //
    task automatic wait_for_config_master_error_position(  );
        begin
            @( config_master_error_position );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_setup_time
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_setup_time>.
    //
    task automatic wait_for_config_setup_time(  );
        begin
            @( config_setup_time );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_hold_time
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_hold_time>.
    //
    task automatic wait_for_config_hold_time(  );
        begin
            @( config_hold_time );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_wr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_wr>.
    //
    task automatic wait_for_config_max_outstanding_wr(  );
        begin
            @( config_max_outstanding_wr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_rd
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_rd>.
    //
    task automatic wait_for_config_max_outstanding_rd(  );
        begin
            @( config_max_outstanding_rd );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_rw
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_rw>.
    //
    task automatic wait_for_config_max_outstanding_rw(  );
        begin
            @( config_max_outstanding_rw );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_is_issuing
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_is_issuing>.
    //
    task automatic wait_for_config_is_issuing(  );
        begin
            @( config_is_issuing );
        end
    endtask


    //-------------------------------------------------------------------------
    // Functions to set global variables with write access
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- set_config_write_ctrl_to_data_mintime
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_write_ctrl_to_data_mintime>.
    //
    // Parameters:
    //     config_write_ctrl_to_data_mintime_param - The value to assign to variable <config_write_ctrl_to_data_mintime>.
    //
    function automatic void set_config_write_ctrl_to_data_mintime( int unsigned config_write_ctrl_to_data_mintime_param );
        config_write_ctrl_to_data_mintime = config_write_ctrl_to_data_mintime_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_master_write_delay
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_master_write_delay>.
    //
    // Parameters:
    //     config_master_write_delay_param - The value to assign to variable <config_master_write_delay>.
    //
    function automatic void set_config_master_write_delay( bit config_master_write_delay_param );
        config_master_write_delay = config_master_write_delay_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_all_assertions
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_enable_all_assertions>.
    //
    // Parameters:
    //     config_enable_all_assertions_param - The value to assign to variable <config_enable_all_assertions>.
    //
    function automatic void set_config_enable_all_assertions( bit config_enable_all_assertions_param );
        config_enable_all_assertions = config_enable_all_assertions_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_assertion
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_enable_assertion>.
    //
    // Parameters:
    //     config_enable_assertion_param - The value to assign to variable <config_enable_assertion>.
    //
    function automatic void set_config_enable_assertion( bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
        config_enable_assertion = config_enable_assertion_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_assertion_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_enable_assertion_param - The value to assign to variable <config_enable_assertion>.
    //
    function automatic void set_config_enable_assertion_index1( int _this_dot_1, bit  config_enable_assertion_param );
        config_enable_assertion[_this_dot_1] = config_enable_assertion_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_start_addr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_slave_start_addr>.
    //
    // Parameters:
    //     config_slave_start_addr_param - The value to assign to variable <config_slave_start_addr>.
    //
    function automatic void set_config_slave_start_addr( bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param );
        config_slave_start_addr = config_slave_start_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_start_addr_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_slave_start_addr_param - The value to assign to variable <config_slave_start_addr>.
    //
    function automatic void set_config_slave_start_addr_index1( int _this_dot_1, bit  config_slave_start_addr_param );
        config_slave_start_addr[_this_dot_1] = config_slave_start_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_end_addr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_slave_end_addr>.
    //
    // Parameters:
    //     config_slave_end_addr_param - The value to assign to variable <config_slave_end_addr>.
    //
    function automatic void set_config_slave_end_addr( bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param );
        config_slave_end_addr = config_slave_end_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_end_addr_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_slave_end_addr_param - The value to assign to variable <config_slave_end_addr>.
    //
    function automatic void set_config_slave_end_addr_index1( int _this_dot_1, bit  config_slave_end_addr_param );
        config_slave_end_addr[_this_dot_1] = config_slave_end_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_support_exclusive_access
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_support_exclusive_access>.
    //
    // Parameters:
    //     config_support_exclusive_access_param - The value to assign to variable <config_support_exclusive_access>.
    //
    function automatic void set_config_support_exclusive_access( bit config_support_exclusive_access_param );
        config_support_exclusive_access = config_support_exclusive_access_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_read_data_reordering_depth
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_read_data_reordering_depth>.
    //
    // Parameters:
    //     config_read_data_reordering_depth_param - The value to assign to variable <config_read_data_reordering_depth>.
    //
    function automatic void set_config_read_data_reordering_depth( int unsigned config_read_data_reordering_depth_param );
        config_read_data_reordering_depth = config_read_data_reordering_depth_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_transaction_time_factor
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_transaction_time_factor>.
    //
    // Parameters:
    //     config_max_transaction_time_factor_param - The value to assign to variable <config_max_transaction_time_factor>.
    //
    function automatic void set_config_max_transaction_time_factor( int unsigned config_max_transaction_time_factor_param );
        config_max_transaction_time_factor = config_max_transaction_time_factor_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_timeout_max_data_transfer
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_timeout_max_data_transfer>.
    //
    // Parameters:
    //     config_timeout_max_data_transfer_param - The value to assign to variable <config_timeout_max_data_transfer>.
    //
    function automatic void set_config_timeout_max_data_transfer( int config_timeout_max_data_transfer_param );
        config_timeout_max_data_transfer = config_timeout_max_data_transfer_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_burst_timeout_factor
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_burst_timeout_factor>.
    //
    // Parameters:
    //     config_burst_timeout_factor_param - The value to assign to variable <config_burst_timeout_factor>.
    //
    function automatic void set_config_burst_timeout_factor( int unsigned config_burst_timeout_factor_param );
        config_burst_timeout_factor = config_burst_timeout_factor_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_AWVALID_assertion_to_AWREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    // Parameters:
    //     config_max_latency_AWVALID_assertion_to_AWREADY_param - The value to assign to variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    function automatic void set_config_max_latency_AWVALID_assertion_to_AWREADY( int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
        config_max_latency_AWVALID_assertion_to_AWREADY = config_max_latency_AWVALID_assertion_to_AWREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_ARVALID_assertion_to_ARREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    // Parameters:
    //     config_max_latency_ARVALID_assertion_to_ARREADY_param - The value to assign to variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    function automatic void set_config_max_latency_ARVALID_assertion_to_ARREADY( int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
        config_max_latency_ARVALID_assertion_to_ARREADY = config_max_latency_ARVALID_assertion_to_ARREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_RVALID_assertion_to_RREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    // Parameters:
    //     config_max_latency_RVALID_assertion_to_RREADY_param - The value to assign to variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    function automatic void set_config_max_latency_RVALID_assertion_to_RREADY( int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
        config_max_latency_RVALID_assertion_to_RREADY = config_max_latency_RVALID_assertion_to_RREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_BVALID_assertion_to_BREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    // Parameters:
    //     config_max_latency_BVALID_assertion_to_BREADY_param - The value to assign to variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    function automatic void set_config_max_latency_BVALID_assertion_to_BREADY( int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
        config_max_latency_BVALID_assertion_to_BREADY = config_max_latency_BVALID_assertion_to_BREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_WVALID_assertion_to_WREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    // Parameters:
    //     config_max_latency_WVALID_assertion_to_WREADY_param - The value to assign to variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    function automatic void set_config_max_latency_WVALID_assertion_to_WREADY( int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
        config_max_latency_WVALID_assertion_to_WREADY = config_max_latency_WVALID_assertion_to_WREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_master_error_position
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_master_error_position>.
    //
    // Parameters:
    //     config_master_error_position_param - The value to assign to variable <config_master_error_position>.
    //
    function automatic void set_config_master_error_position( axi_error_e config_master_error_position_param );
        config_master_error_position = config_master_error_position_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_setup_time
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_setup_time>.
    //
    // Parameters:
    //     config_setup_time_param - The value to assign to variable <config_setup_time>.
    //
    function automatic void set_config_setup_time( int config_setup_time_param );
        config_setup_time = config_setup_time_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_hold_time
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_hold_time>.
    //
    // Parameters:
    //     config_hold_time_param - The value to assign to variable <config_hold_time>.
    //
    function automatic void set_config_hold_time( int config_hold_time_param );
        config_hold_time = config_hold_time_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_wr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_wr>.
    //
    // Parameters:
    //     config_max_outstanding_wr_param - The value to assign to variable <config_max_outstanding_wr>.
    //
    function automatic void set_config_max_outstanding_wr( int config_max_outstanding_wr_param );
        config_max_outstanding_wr = config_max_outstanding_wr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_rd
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_rd>.
    //
    // Parameters:
    //     config_max_outstanding_rd_param - The value to assign to variable <config_max_outstanding_rd>.
    //
    function automatic void set_config_max_outstanding_rd( int config_max_outstanding_rd_param );
        config_max_outstanding_rd = config_max_outstanding_rd_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_rw
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_rw>.
    //
    // Parameters:
    //     config_max_outstanding_rw_param - The value to assign to variable <config_max_outstanding_rw>.
    //
    function automatic void set_config_max_outstanding_rw( int config_max_outstanding_rw_param );
        config_max_outstanding_rw = config_max_outstanding_rw_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_is_issuing
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_is_issuing>.
    //
    // Parameters:
    //     config_is_issuing_param - The value to assign to variable <config_is_issuing>.
    //
    function automatic void set_config_is_issuing( bit config_is_issuing_param );
        config_is_issuing = config_is_issuing_param;
    endfunction


    //-------------------------------------------------------------------------
    // Functions to get global variables with read access
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- get_config_write_ctrl_to_data_mintime
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_write_ctrl_to_data_mintime>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_write_ctrl_to_data_mintime>.
    //
    function automatic int unsigned get_config_write_ctrl_to_data_mintime(  );
        return config_write_ctrl_to_data_mintime;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_master_write_delay
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_master_write_delay>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_master_write_delay>.
    //
    function automatic bit get_config_master_write_delay(  );
        axi_get_deprecated_config_master_write_delay_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_master_write_delay;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_all_assertions
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_enable_all_assertions>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_enable_all_assertions>.
    //
    function automatic bit get_config_enable_all_assertions(  );
        return config_enable_all_assertions;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_assertion
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_enable_assertion>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_enable_assertion>.
    //
    function automatic bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]   get_config_enable_assertion(  );
        return config_enable_assertion;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_assertion_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_enable_assertion>.
    //
    function automatic bit   get_config_enable_assertion_index1( int _this_dot_1 );
        return config_enable_assertion[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_start_addr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_slave_start_addr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_slave_start_addr>.
    //
    function automatic bit [((AXI_ADDRESS_WIDTH) - 1):0]   get_config_slave_start_addr(  );
        axi_get_deprecated_config_slave_start_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_start_addr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_start_addr_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_slave_start_addr>.
    //
    function automatic bit   get_config_slave_start_addr_index1( int _this_dot_1 );
        axi_get_deprecated_config_slave_start_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_start_addr[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_end_addr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_slave_end_addr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_slave_end_addr>.
    //
    function automatic bit [((AXI_ADDRESS_WIDTH) - 1):0]   get_config_slave_end_addr(  );
        axi_get_deprecated_config_slave_end_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_end_addr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_end_addr_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_slave_end_addr>.
    //
    function automatic bit   get_config_slave_end_addr_index1( int _this_dot_1 );
        axi_get_deprecated_config_slave_end_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_end_addr[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_support_exclusive_access
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_support_exclusive_access>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_support_exclusive_access>.
    //
    function automatic bit get_config_support_exclusive_access(  );
        return config_support_exclusive_access;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_read_data_reordering_depth
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_read_data_reordering_depth>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_read_data_reordering_depth>.
    //
    function automatic int unsigned get_config_read_data_reordering_depth(  );
        return config_read_data_reordering_depth;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_transaction_time_factor
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_transaction_time_factor>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_transaction_time_factor>.
    //
    function automatic int unsigned get_config_max_transaction_time_factor(  );
        return config_max_transaction_time_factor;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_timeout_max_data_transfer
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_timeout_max_data_transfer>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_timeout_max_data_transfer>.
    //
    function automatic int get_config_timeout_max_data_transfer(  );
        return config_timeout_max_data_transfer;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_burst_timeout_factor
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_burst_timeout_factor>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_burst_timeout_factor>.
    //
    function automatic int unsigned get_config_burst_timeout_factor(  );
        return config_burst_timeout_factor;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_AWVALID_assertion_to_AWREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    function automatic int unsigned get_config_max_latency_AWVALID_assertion_to_AWREADY(  );
        return config_max_latency_AWVALID_assertion_to_AWREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_ARVALID_assertion_to_ARREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    function automatic int unsigned get_config_max_latency_ARVALID_assertion_to_ARREADY(  );
        return config_max_latency_ARVALID_assertion_to_ARREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_RVALID_assertion_to_RREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    function automatic int unsigned get_config_max_latency_RVALID_assertion_to_RREADY(  );
        return config_max_latency_RVALID_assertion_to_RREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_BVALID_assertion_to_BREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    function automatic int unsigned get_config_max_latency_BVALID_assertion_to_BREADY(  );
        return config_max_latency_BVALID_assertion_to_BREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_WVALID_assertion_to_WREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    function automatic int unsigned get_config_max_latency_WVALID_assertion_to_WREADY(  );
        return config_max_latency_WVALID_assertion_to_WREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_master_error_position
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_master_error_position>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_master_error_position>.
    //
    function automatic axi_error_e get_config_master_error_position(  );
        axi_get_deprecated_config_master_error_position_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_master_error_position;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_setup_time
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_setup_time>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_setup_time>.
    //
    function automatic int get_config_setup_time(  );
        return config_setup_time;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_hold_time
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_hold_time>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_hold_time>.
    //
    function automatic int get_config_hold_time(  );
        return config_hold_time;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_wr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_wr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_wr>.
    //
    function automatic int get_config_max_outstanding_wr(  );
        return config_max_outstanding_wr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_rd
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_rd>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_rd>.
    //
    function automatic int get_config_max_outstanding_rd(  );
        return config_max_outstanding_rd;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_rw
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_rw>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_rw>.
    //
    function automatic int get_config_max_outstanding_rw(  );
        return config_max_outstanding_rw;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_is_issuing
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_is_issuing>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_is_issuing>.
    //
    function automatic bit get_config_is_issuing(  );
        return config_is_issuing;
    endfunction


    //-------------------------------------------------------------------------
    // Functions to set/get generic interface configuration
    //-------------------------------------------------------------------------

    function void set_interface
    (
        input int what = 0,
        input int arg1 = 0,
        input int arg2 = 0,
        input int arg3 = 0,
        input int arg4 = 0,
        input int arg5 = 0,
        input int arg6 = 0,
        input int arg7 = 0,
        input int arg8 = 0,
        input int arg9 = 0,
        input int arg10 = 0
    );
        axi_set_interface( what, arg1, arg2, arg3, arg4, arg5, arg6, arg7, arg8, arg9, arg10 );
    endfunction

    function int get_interface
    (
        input int what = 0,
        input int arg1 = 0,
        input int arg2 = 0,
        input int arg3 = 0,
        input int arg4 = 0,
        input int arg5 = 0,
        input int arg6 = 0,
        input int arg7 = 0,
        input int arg8 = 0,
        input int arg9 = 0
    );
        return axi_get_interface( what, arg1, arg2, arg3, arg4, arg5, arg6, arg7, arg8, arg9 );
    endfunction

    //-------------------------------------------------------------------------
    // Functions to get the hierarchic name of this interface
    //-------------------------------------------------------------------------
    function string get_full_name();
        return axi_get_full_name();
    endfunction

    //--------------------------------------------------------------------------
    //
    // Group:- Monitor Value Change on Variable
    //
    //--------------------------------------------------------------------------

    function automatic void axi_local_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( ref int unsigned config_write_ctrl_to_data_mintime_param );
            axi_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( _interface_ref,config_write_ctrl_to_data_mintime); // DPI call to imported task
        
            axi_propagate_config_write_ctrl_to_data_mintime_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( config_write_ctrl_to_data_mintime );
            end
        end
    end

    function automatic void axi_local_set_config_master_write_delay_from_SystemVerilog( ref bit config_master_write_delay_param );
            axi_set_config_master_write_delay_from_SystemVerilog( _interface_ref,config_master_write_delay); // DPI call to imported task
        
            axi_propagate_config_master_write_delay_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_master_write_delay_from_SystemVerilog( config_master_write_delay );
            end
        end
    end

    function automatic void axi_local_set_config_enable_all_assertions_from_SystemVerilog( ref bit config_enable_all_assertions_param );
            axi_set_config_enable_all_assertions_from_SystemVerilog( _interface_ref,config_enable_all_assertions); // DPI call to imported task
        
            axi_propagate_config_enable_all_assertions_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_enable_all_assertions_from_SystemVerilog( config_enable_all_assertions );
            end
        end
    end

    function automatic void axi_local_set_config_enable_assertion_from_SystemVerilog( ref bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
            axi_set_config_enable_assertion_from_SystemVerilog( _interface_ref,config_enable_assertion); // DPI call to imported task
        
            axi_propagate_config_enable_assertion_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_enable_assertion_from_SystemVerilog( config_enable_assertion );
            end
        end
    end

    function automatic void axi_local_set_config_slave_start_addr_from_SystemVerilog( ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ADDRESS_WIDTH ); _this_dot_1++)
        begin
            axi_set_config_slave_start_addr_from_SystemVerilog_index1( _interface_ref,_this_dot_1,config_slave_start_addr[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
            axi_propagate_config_slave_start_addr_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_slave_start_addr_from_SystemVerilog( config_slave_start_addr );
            end
        end
    end

    function automatic void axi_local_set_config_slave_end_addr_from_SystemVerilog( ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ADDRESS_WIDTH ); _this_dot_1++)
        begin
            axi_set_config_slave_end_addr_from_SystemVerilog_index1( _interface_ref,_this_dot_1,config_slave_end_addr[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
            axi_propagate_config_slave_end_addr_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_slave_end_addr_from_SystemVerilog( config_slave_end_addr );
            end
        end
    end

    function automatic void axi_local_set_config_support_exclusive_access_from_SystemVerilog( ref bit config_support_exclusive_access_param );
            axi_set_config_support_exclusive_access_from_SystemVerilog( _interface_ref,config_support_exclusive_access); // DPI call to imported task
        
            axi_propagate_config_support_exclusive_access_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_support_exclusive_access_from_SystemVerilog( config_support_exclusive_access );
            end
        end
    end

    function automatic void axi_local_set_config_read_data_reordering_depth_from_SystemVerilog( ref int unsigned config_read_data_reordering_depth_param );
            axi_set_config_read_data_reordering_depth_from_SystemVerilog( _interface_ref,config_read_data_reordering_depth); // DPI call to imported task
        
            axi_propagate_config_read_data_reordering_depth_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_read_data_reordering_depth_from_SystemVerilog( config_read_data_reordering_depth );
            end
        end
    end

    function automatic void axi_local_set_config_max_transaction_time_factor_from_SystemVerilog( ref int unsigned config_max_transaction_time_factor_param );
            axi_set_config_max_transaction_time_factor_from_SystemVerilog( _interface_ref,config_max_transaction_time_factor); // DPI call to imported task
        
            axi_propagate_config_max_transaction_time_factor_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_transaction_time_factor_from_SystemVerilog( config_max_transaction_time_factor );
            end
        end
    end

    function automatic void axi_local_set_config_timeout_max_data_transfer_from_SystemVerilog( ref int config_timeout_max_data_transfer_param );
            axi_set_config_timeout_max_data_transfer_from_SystemVerilog( _interface_ref,config_timeout_max_data_transfer); // DPI call to imported task
        
            axi_propagate_config_timeout_max_data_transfer_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_timeout_max_data_transfer_from_SystemVerilog( config_timeout_max_data_transfer );
            end
        end
    end

    function automatic void axi_local_set_config_burst_timeout_factor_from_SystemVerilog( ref int unsigned config_burst_timeout_factor_param );
            axi_set_config_burst_timeout_factor_from_SystemVerilog( _interface_ref,config_burst_timeout_factor); // DPI call to imported task
        
            axi_propagate_config_burst_timeout_factor_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_burst_timeout_factor_from_SystemVerilog( config_burst_timeout_factor );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( ref int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
            axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( _interface_ref,config_max_latency_AWVALID_assertion_to_AWREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( config_max_latency_AWVALID_assertion_to_AWREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( ref int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
            axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( _interface_ref,config_max_latency_ARVALID_assertion_to_ARREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( config_max_latency_ARVALID_assertion_to_ARREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( ref int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
            axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( _interface_ref,config_max_latency_RVALID_assertion_to_RREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( config_max_latency_RVALID_assertion_to_RREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( ref int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
            axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( _interface_ref,config_max_latency_BVALID_assertion_to_BREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( config_max_latency_BVALID_assertion_to_BREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( ref int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
            axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( _interface_ref,config_max_latency_WVALID_assertion_to_WREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( config_max_latency_WVALID_assertion_to_WREADY );
            end
        end
    end

    function automatic void axi_local_set_config_master_error_position_from_SystemVerilog( ref axi_error_e config_master_error_position_param );
            axi_set_config_master_error_position_from_SystemVerilog( _interface_ref,config_master_error_position); // DPI call to imported task
        
            axi_propagate_config_master_error_position_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_master_error_position_from_SystemVerilog( config_master_error_position );
            end
        end
    end

    function automatic void axi_local_set_config_setup_time_from_SystemVerilog( ref int config_setup_time_param );
            axi_set_config_setup_time_from_SystemVerilog( _interface_ref,config_setup_time); // DPI call to imported task
        
            axi_propagate_config_setup_time_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_setup_time_from_SystemVerilog( config_setup_time );
            end
        end
    end

    function automatic void axi_local_set_config_hold_time_from_SystemVerilog( ref int config_hold_time_param );
            axi_set_config_hold_time_from_SystemVerilog( _interface_ref,config_hold_time); // DPI call to imported task
        
            axi_propagate_config_hold_time_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_hold_time_from_SystemVerilog( config_hold_time );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_wr_from_SystemVerilog( ref int config_max_outstanding_wr_param );
            axi_set_config_max_outstanding_wr_from_SystemVerilog( _interface_ref,config_max_outstanding_wr); // DPI call to imported task
        
            axi_propagate_config_max_outstanding_wr_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_wr_from_SystemVerilog( config_max_outstanding_wr );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_rd_from_SystemVerilog( ref int config_max_outstanding_rd_param );
            axi_set_config_max_outstanding_rd_from_SystemVerilog( _interface_ref,config_max_outstanding_rd); // DPI call to imported task
        
            axi_propagate_config_max_outstanding_rd_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_rd_from_SystemVerilog( config_max_outstanding_rd );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_rw_from_SystemVerilog( ref int config_max_outstanding_rw_param );
            axi_set_config_max_outstanding_rw_from_SystemVerilog( _interface_ref,config_max_outstanding_rw); // DPI call to imported task
        
            axi_propagate_config_max_outstanding_rw_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_rw_from_SystemVerilog( config_max_outstanding_rw );
            end
        end
    end

    function automatic void axi_local_set_config_is_issuing_from_SystemVerilog( ref bit config_is_issuing_param );
            axi_set_config_is_issuing_from_SystemVerilog( _interface_ref,config_is_issuing); // DPI call to imported task
        
            axi_propagate_config_is_issuing_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_is_issuing_from_SystemVerilog( config_is_issuing );
            end
        end
    end

    //-------------------------------------------------------------------------
    // Transaction interface
    //-------------------------------------------------------------------------

    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_rw_transaction_addr;
    function void axi_get_temp_static_rw_transaction_addr( input int _d1, output bit  _value );
        _value = temp_static_rw_transaction_addr[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_addr( input int _d1, input bit  _value );
        temp_static_rw_transaction_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_rw_transaction_id;
    function void axi_get_temp_static_rw_transaction_id( input int _d1, output bit  _value );
        _value = temp_static_rw_transaction_id[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_id( input int _d1, input bit  _value );
        temp_static_rw_transaction_id[_d1] = _value;
    endfunction
    bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] temp_static_rw_transaction_data_words [];
    function void axi_get_temp_static_rw_transaction_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_rw_transaction_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_rw_transaction_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_rw_transaction_data_words[_d1][_d2] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] temp_static_rw_transaction_write_strobes [];
    function void axi_get_temp_static_rw_transaction_write_strobes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_rw_transaction_write_strobes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_rw_transaction_write_strobes( input int _d1, input int _d2, input bit _value );
        temp_static_rw_transaction_write_strobes[_d1][_d2] = _value;
    endfunction
    axi_response_e temp_static_rw_transaction_resp[];
    function void axi_get_temp_static_rw_transaction_resp( input int _d1, output axi_response_e _value );
        _value = temp_static_rw_transaction_resp[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_resp( input int _d1, input axi_response_e _value );
        temp_static_rw_transaction_resp[_d1] = _value;
    endfunction
    bit [7:0] temp_static_rw_transaction_data_user [];
    function void axi_get_temp_static_rw_transaction_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_rw_transaction_data_user[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_rw_transaction_data_user[_d1] = _value;
    endfunction
    int temp_static_rw_transaction_write_data_beats_delay[];
    function void axi_get_temp_static_rw_transaction_write_data_beats_delay( input int _d1, output int _value );
        _value = temp_static_rw_transaction_write_data_beats_delay[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_write_data_beats_delay( input int _d1, input int _value );
        temp_static_rw_transaction_write_data_beats_delay[_d1] = _value;
    endfunction
    int temp_static_rw_transaction_data_valid_delay[];
    function void axi_get_temp_static_rw_transaction_data_valid_delay( input int _d1, output int _value );
        _value = temp_static_rw_transaction_data_valid_delay[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_data_valid_delay( input int _d1, input int _value );
        temp_static_rw_transaction_data_valid_delay[_d1] = _value;
    endfunction
    int temp_static_rw_transaction_data_ready_delay[];
    function void axi_get_temp_static_rw_transaction_data_ready_delay( input int _d1, output int _value );
        _value = temp_static_rw_transaction_data_ready_delay[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_data_ready_delay( input int _d1, input int _value );
        temp_static_rw_transaction_data_ready_delay[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_AXI_read_addr;
    function void axi_get_temp_static_AXI_read_addr( input int _d1, output bit  _value );
        _value = temp_static_AXI_read_addr[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_addr( input int _d1, input bit  _value );
        temp_static_AXI_read_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_AXI_read_id;
    function void axi_get_temp_static_AXI_read_id( input int _d1, output bit  _value );
        _value = temp_static_AXI_read_id[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_id( input int _d1, input bit  _value );
        temp_static_AXI_read_id[_d1] = _value;
    endfunction
    bit [((AXI_RDATA_WIDTH) - 1):0] temp_static_AXI_read_data_words [];
    function void axi_get_temp_static_AXI_read_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_AXI_read_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_AXI_read_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_AXI_read_data_words[_d1][_d2] = _value;
    endfunction
    axi_response_e temp_static_AXI_read_resp[];
    function void axi_get_temp_static_AXI_read_resp( input int _d1, output axi_response_e _value );
        _value = temp_static_AXI_read_resp[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_resp( input int _d1, input axi_response_e _value );
        temp_static_AXI_read_resp[_d1] = _value;
    endfunction
    bit [7:0] temp_static_AXI_read_data_user [];
    function void axi_get_temp_static_AXI_read_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_AXI_read_data_user[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_AXI_read_data_user[_d1] = _value;
    endfunction
    longint temp_static_AXI_read_data_start_time[];
    function void axi_get_temp_static_AXI_read_data_start_time( input int _d1, output longint _value );
        _value = temp_static_AXI_read_data_start_time[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_data_start_time( input int _d1, input longint _value );
        temp_static_AXI_read_data_start_time[_d1] = _value;
    endfunction
    longint temp_static_AXI_read_data_end_time[];
    function void axi_get_temp_static_AXI_read_data_end_time( input int _d1, output longint _value );
        _value = temp_static_AXI_read_data_end_time[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_data_end_time( input int _d1, input longint _value );
        temp_static_AXI_read_data_end_time[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_AXI_write_addr;
    function void axi_get_temp_static_AXI_write_addr( input int _d1, output bit  _value );
        _value = temp_static_AXI_write_addr[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_addr( input int _d1, input bit  _value );
        temp_static_AXI_write_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_AXI_write_id;
    function void axi_get_temp_static_AXI_write_id( input int _d1, output bit  _value );
        _value = temp_static_AXI_write_id[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_id( input int _d1, input bit  _value );
        temp_static_AXI_write_id[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0] temp_static_AXI_write_data_words [];
    function void axi_get_temp_static_AXI_write_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_AXI_write_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_AXI_write_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_AXI_write_data_words[_d1][_d2] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] temp_static_AXI_write_write_strobes [];
    function void axi_get_temp_static_AXI_write_write_strobes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_AXI_write_write_strobes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_AXI_write_write_strobes( input int _d1, input int _d2, input bit _value );
        temp_static_AXI_write_write_strobes[_d1][_d2] = _value;
    endfunction
    bit [7:0] temp_static_AXI_write_data_user [];
    function void axi_get_temp_static_AXI_write_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_AXI_write_data_user[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_AXI_write_data_user[_d1] = _value;
    endfunction
    int temp_static_AXI_write_write_data_beats_delay[];
    function void axi_get_temp_static_AXI_write_write_data_beats_delay( input int _d1, output int _value );
        _value = temp_static_AXI_write_write_data_beats_delay[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_write_data_beats_delay( input int _d1, input int _value );
        temp_static_AXI_write_write_data_beats_delay[_d1] = _value;
    endfunction
    longint temp_static_AXI_write_data_start_time[];
    function void axi_get_temp_static_AXI_write_data_start_time( input int _d1, output longint _value );
        _value = temp_static_AXI_write_data_start_time[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_data_start_time( input int _d1, input longint _value );
        temp_static_AXI_write_data_start_time[_d1] = _value;
    endfunction
    longint temp_static_AXI_write_data_end_time[];
    function void axi_get_temp_static_AXI_write_data_end_time( input int _d1, output longint _value );
        _value = temp_static_AXI_write_data_end_time[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_data_end_time( input int _d1, input longint _value );
        temp_static_AXI_write_data_end_time[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0] temp_static_data_resp_data_words [];
    function void axi_get_temp_static_data_resp_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_data_resp_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_data_resp_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_data_resp_data_words[_d1][_d2] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] temp_static_data_resp_write_strobes [];
    function void axi_get_temp_static_data_resp_write_strobes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_data_resp_write_strobes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_data_resp_write_strobes( input int _d1, input int _d2, input bit _value );
        temp_static_data_resp_write_strobes[_d1][_d2] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_data_resp_id;
    function void axi_get_temp_static_data_resp_id( input int _d1, output bit  _value );
        _value = temp_static_data_resp_id[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_id( input int _d1, input bit  _value );
        temp_static_data_resp_id[_d1] = _value;
    endfunction
    bit [7:0] temp_static_data_resp_data_user [];
    function void axi_get_temp_static_data_resp_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_data_resp_data_user[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_data_resp_data_user[_d1] = _value;
    endfunction
    int temp_static_data_resp_write_data_beats_delay[];
    function void axi_get_temp_static_data_resp_write_data_beats_delay( input int _d1, output int _value );
        _value = temp_static_data_resp_write_data_beats_delay[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_write_data_beats_delay( input int _d1, input int _value );
        temp_static_data_resp_write_data_beats_delay[_d1] = _value;
    endfunction
    longint temp_static_data_resp_data_beat_start_time[];
    function void axi_get_temp_static_data_resp_data_beat_start_time( input int _d1, output longint _value );
        _value = temp_static_data_resp_data_beat_start_time[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_data_beat_start_time( input int _d1, input longint _value );
        temp_static_data_resp_data_beat_start_time[_d1] = _value;
    endfunction
    longint temp_static_data_resp_data_beat_end_time[];
    function void axi_get_temp_static_data_resp_data_beat_end_time( input int _d1, output longint _value );
        _value = temp_static_data_resp_data_beat_end_time[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_data_beat_end_time( input int _d1, input longint _value );
        temp_static_data_resp_data_beat_end_time[_d1] = _value;
    endfunction
    bit [((AXI_RDATA_WIDTH) - 1):0] temp_static_read_data_burst_data_words [];
    function void axi_get_temp_static_read_data_burst_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_read_data_burst_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_read_data_burst_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_read_data_burst_data_words[_d1][_d2] = _value;
    endfunction
    axi_response_e temp_static_read_data_burst_resp[];
    function void axi_get_temp_static_read_data_burst_resp( input int _d1, output axi_response_e _value );
        _value = temp_static_read_data_burst_resp[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_resp( input int _d1, input axi_response_e _value );
        temp_static_read_data_burst_resp[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_data_burst_id;
    function void axi_get_temp_static_read_data_burst_id( input int _d1, output bit  _value );
        _value = temp_static_read_data_burst_id[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_id( input int _d1, input bit  _value );
        temp_static_read_data_burst_id[_d1] = _value;
    endfunction
    bit [7:0] temp_static_read_data_burst_data_user [];
    function void axi_get_temp_static_read_data_burst_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_read_data_burst_data_user[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_read_data_burst_data_user[_d1] = _value;
    endfunction
    longint temp_static_read_data_burst_data_start_time[];
    function void axi_get_temp_static_read_data_burst_data_start_time( input int _d1, output longint _value );
        _value = temp_static_read_data_burst_data_start_time[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_data_start_time( input int _d1, input longint _value );
        temp_static_read_data_burst_data_start_time[_d1] = _value;
    endfunction
    longint temp_static_read_data_burst_data_end_time[];
    function void axi_get_temp_static_read_data_burst_data_end_time( input int _d1, output longint _value );
        _value = temp_static_read_data_burst_data_end_time[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_data_end_time( input int _d1, input longint _value );
        temp_static_read_data_burst_data_end_time[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0] temp_static_write_data_burst_data_words [];
    function void axi_get_temp_static_write_data_burst_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_write_data_burst_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_write_data_burst_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_write_data_burst_data_words[_d1][_d2] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] temp_static_write_data_burst_write_strobes [];
    function void axi_get_temp_static_write_data_burst_write_strobes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_write_data_burst_write_strobes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_write_data_burst_write_strobes( input int _d1, input int _d2, input bit _value );
        temp_static_write_data_burst_write_strobes[_d1][_d2] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_data_burst_id;
    function void axi_get_temp_static_write_data_burst_id( input int _d1, output bit  _value );
        _value = temp_static_write_data_burst_id[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_id( input int _d1, input bit  _value );
        temp_static_write_data_burst_id[_d1] = _value;
    endfunction
    bit [7:0] temp_static_write_data_burst_data_user [];
    function void axi_get_temp_static_write_data_burst_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_write_data_burst_data_user[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_write_data_burst_data_user[_d1] = _value;
    endfunction
    int temp_static_write_data_burst_write_data_beats_delay[];
    function void axi_get_temp_static_write_data_burst_write_data_beats_delay( input int _d1, output int _value );
        _value = temp_static_write_data_burst_write_data_beats_delay[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_write_data_beats_delay( input int _d1, input int _value );
        temp_static_write_data_burst_write_data_beats_delay[_d1] = _value;
    endfunction
    longint temp_static_write_data_burst_data_start_time[];
    function void axi_get_temp_static_write_data_burst_data_start_time( input int _d1, output longint _value );
        _value = temp_static_write_data_burst_data_start_time[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_data_start_time( input int _d1, input longint _value );
        temp_static_write_data_burst_data_start_time[_d1] = _value;
    endfunction
    longint temp_static_write_data_burst_data_end_time[];
    function void axi_get_temp_static_write_data_burst_data_end_time( input int _d1, output longint _value );
        _value = temp_static_write_data_burst_data_end_time[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_data_end_time( input int _d1, input longint _value );
        temp_static_write_data_burst_data_end_time[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_read_addr_channel_phase_addr;
    function void axi_get_temp_static_read_addr_channel_phase_addr( input int _d1, output bit  _value );
        _value = temp_static_read_addr_channel_phase_addr[_d1];
    endfunction
    function void axi_set_temp_static_read_addr_channel_phase_addr( input int _d1, input bit  _value );
        temp_static_read_addr_channel_phase_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_addr_channel_phase_id;
    function void axi_get_temp_static_read_addr_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_read_addr_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_read_addr_channel_phase_id( input int _d1, input bit  _value );
        temp_static_read_addr_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_RDATA_WIDTH) - 1):0]  temp_static_read_channel_phase_data;
    function void axi_get_temp_static_read_channel_phase_data( input int _d1, output bit  _value );
        _value = temp_static_read_channel_phase_data[_d1];
    endfunction
    function void axi_set_temp_static_read_channel_phase_data( input int _d1, input bit  _value );
        temp_static_read_channel_phase_data[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_channel_phase_id;
    function void axi_get_temp_static_read_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_read_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_read_channel_phase_id( input int _d1, input bit  _value );
        temp_static_read_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_write_addr_channel_phase_addr;
    function void axi_get_temp_static_write_addr_channel_phase_addr( input int _d1, output bit  _value );
        _value = temp_static_write_addr_channel_phase_addr[_d1];
    endfunction
    function void axi_set_temp_static_write_addr_channel_phase_addr( input int _d1, input bit  _value );
        temp_static_write_addr_channel_phase_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_addr_channel_phase_id;
    function void axi_get_temp_static_write_addr_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_write_addr_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_write_addr_channel_phase_id( input int _d1, input bit  _value );
        temp_static_write_addr_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0]  temp_static_write_channel_phase_data;
    function void axi_get_temp_static_write_channel_phase_data( input int _d1, output bit  _value );
        _value = temp_static_write_channel_phase_data[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_phase_data( input int _d1, input bit  _value );
        temp_static_write_channel_phase_data[_d1] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  temp_static_write_channel_phase_write_strobes;
    function void axi_get_temp_static_write_channel_phase_write_strobes( input int _d1, output bit  _value );
        _value = temp_static_write_channel_phase_write_strobes[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_phase_write_strobes( input int _d1, input bit  _value );
        temp_static_write_channel_phase_write_strobes[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_channel_phase_id;
    function void axi_get_temp_static_write_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_write_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_phase_id( input int _d1, input bit  _value );
        temp_static_write_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_resp_channel_phase_id;
    function void axi_get_temp_static_write_resp_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_write_resp_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_write_resp_channel_phase_id( input int _d1, input bit  _value );
        temp_static_write_resp_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_read_addr_channel_cycle_addr;
    function void axi_get_temp_static_read_addr_channel_cycle_addr( input int _d1, output bit  _value );
        _value = temp_static_read_addr_channel_cycle_addr[_d1];
    endfunction
    function void axi_set_temp_static_read_addr_channel_cycle_addr( input int _d1, input bit  _value );
        temp_static_read_addr_channel_cycle_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_addr_channel_cycle_id;
    function void axi_get_temp_static_read_addr_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_read_addr_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_read_addr_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_read_addr_channel_cycle_id[_d1] = _value;
    endfunction
    bit [((AXI_RDATA_WIDTH) - 1):0]  temp_static_read_channel_cycle_data;
    function void axi_get_temp_static_read_channel_cycle_data( input int _d1, output bit  _value );
        _value = temp_static_read_channel_cycle_data[_d1];
    endfunction
    function void axi_set_temp_static_read_channel_cycle_data( input int _d1, input bit  _value );
        temp_static_read_channel_cycle_data[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_channel_cycle_id;
    function void axi_get_temp_static_read_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_read_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_read_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_read_channel_cycle_id[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_write_addr_channel_cycle_addr;
    function void axi_get_temp_static_write_addr_channel_cycle_addr( input int _d1, output bit  _value );
        _value = temp_static_write_addr_channel_cycle_addr[_d1];
    endfunction
    function void axi_set_temp_static_write_addr_channel_cycle_addr( input int _d1, input bit  _value );
        temp_static_write_addr_channel_cycle_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_addr_channel_cycle_id;
    function void axi_get_temp_static_write_addr_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_write_addr_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_write_addr_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_write_addr_channel_cycle_id[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0]  temp_static_write_channel_cycle_data;
    function void axi_get_temp_static_write_channel_cycle_data( input int _d1, output bit  _value );
        _value = temp_static_write_channel_cycle_data[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_cycle_data( input int _d1, input bit  _value );
        temp_static_write_channel_cycle_data[_d1] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  temp_static_write_channel_cycle_strb;
    function void axi_get_temp_static_write_channel_cycle_strb( input int _d1, output bit  _value );
        _value = temp_static_write_channel_cycle_strb[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_cycle_strb( input int _d1, input bit  _value );
        temp_static_write_channel_cycle_strb[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_channel_cycle_id;
    function void axi_get_temp_static_write_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_write_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_write_channel_cycle_id[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_resp_channel_cycle_id;
    function void axi_get_temp_static_write_resp_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_write_resp_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_write_resp_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_write_resp_channel_cycle_id[_d1] = _value;
    endfunction
    task automatic dvc_activate_rw_transaction
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp[],
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref axi_rw_e read_or_write,
        ref int address_to_data_latency,
        ref int data_to_response_latency,
        ref int write_address_to_data_delay,
        ref int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        ref int address_valid_delay,
        ref int data_valid_delay[],
        ref int write_response_valid_delay,
        ref int address_ready_delay,
        ref int data_ready_delay[],
        ref int write_response_ready_delay,
        ref bit write_data_with_address,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_valid_delay_DIMS0;
                automatic int data_ready_delay_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_rw_transaction_addr = addr;
            temp_static_rw_transaction_id = id;
            data_words_DIMS0 = data_words.size();
            temp_static_rw_transaction_data_words = data_words;
            write_strobes_DIMS0 = write_strobes.size();
            temp_static_rw_transaction_write_strobes = write_strobes;
            resp_DIMS0 = resp.size();
            temp_static_rw_transaction_resp = resp;
            data_user_DIMS0 = data_user.size();
            temp_static_rw_transaction_data_user = data_user;
            write_data_beats_delay_DIMS0 = write_data_beats_delay.size();
            temp_static_rw_transaction_write_data_beats_delay = write_data_beats_delay;
            data_valid_delay_DIMS0 = data_valid_delay.size();
            temp_static_rw_transaction_data_valid_delay = data_valid_delay;
            data_ready_delay_DIMS0 = data_ready_delay.size();
            temp_static_rw_transaction_data_ready_delay = data_ready_delay;
            // Call function to provide sized params and ingoing unsized params sizes.
            // In addition gets back updated sizes of unsized params.
            axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, data_words_DIMS0, write_strobes_DIMS0, resp_DIMS0, addr_user, data_user_DIMS0, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay_DIMS0, address_valid_delay, data_valid_delay_DIMS0, write_response_valid_delay, address_ready_delay, data_ready_delay_DIMS0, write_response_ready_delay, write_data_with_address, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_rw_transaction_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_write_strobes.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_rw_transaction_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_write_data_beats_delay.delete();
            end
            if (data_valid_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_valid_delay = new [data_valid_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_valid_delay.delete();
            end
            if (data_ready_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_ready_delay = new [data_ready_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_ready_delay.delete();
            end
            // Call function to get the sized params
            axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, addr_user, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, address_valid_delay, write_response_valid_delay, address_ready_delay, write_response_ready_delay, write_data_with_address, _unit_id); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_rw_transaction_addr;
            id = temp_static_rw_transaction_id;
            data_words = temp_static_rw_transaction_data_words;
            temp_static_rw_transaction_data_words.delete();
            write_strobes = temp_static_rw_transaction_write_strobes;
            temp_static_rw_transaction_write_strobes.delete();
            resp = temp_static_rw_transaction_resp;
            temp_static_rw_transaction_resp.delete();
            data_user = temp_static_rw_transaction_data_user;
            temp_static_rw_transaction_data_user.delete();
            write_data_beats_delay = temp_static_rw_transaction_write_data_beats_delay;
            temp_static_rw_transaction_write_data_beats_delay.delete();
            data_valid_delay = temp_static_rw_transaction_data_valid_delay;
            temp_static_rw_transaction_data_valid_delay.delete();
            data_ready_delay = temp_static_rw_transaction_data_ready_delay;
            temp_static_rw_transaction_data_ready_delay.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_rw_transaction
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp[],
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output axi_rw_e read_or_write,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        output int address_valid_delay,
        ref int data_valid_delay[],
        output int write_response_valid_delay,
        output int address_ready_delay,
        ref int data_ready_delay[],
        output int write_response_ready_delay,
        output bit write_data_with_address,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_valid_delay_DIMS0;
                automatic int data_ready_delay_DIMS0;
            // Call function to get unsized params sizes.
            axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, resp_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_valid_delay_DIMS0, data_ready_delay_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_rw_transaction_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_write_strobes.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_rw_transaction_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_write_data_beats_delay.delete();
            end
            if (data_valid_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_valid_delay = new [data_valid_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_valid_delay.delete();
            end
            if (data_ready_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_ready_delay = new [data_ready_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_ready_delay.delete();
            end
            // Call function to get the sized params
            axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, addr_user, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, address_valid_delay, write_response_valid_delay, address_ready_delay, write_response_ready_delay, write_data_with_address, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_rw_transaction_addr;
            id = temp_static_rw_transaction_id;
            data_words = temp_static_rw_transaction_data_words;
            temp_static_rw_transaction_data_words.delete();
            write_strobes = temp_static_rw_transaction_write_strobes;
            temp_static_rw_transaction_write_strobes.delete();
            resp = temp_static_rw_transaction_resp;
            temp_static_rw_transaction_resp.delete();
            data_user = temp_static_rw_transaction_data_user;
            temp_static_rw_transaction_data_user.delete();
            write_data_beats_delay = temp_static_rw_transaction_write_data_beats_delay;
            temp_static_rw_transaction_write_data_beats_delay.delete();
            data_valid_delay = temp_static_rw_transaction_data_valid_delay;
            temp_static_rw_transaction_data_valid_delay.delete();
            data_ready_delay = temp_static_rw_transaction_data_ready_delay;
            temp_static_rw_transaction_data_ready_delay.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_AXI_read
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref int address_to_data_latency,
        ref longint addr_start_time,
        ref longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        ref int address_valid_delay,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_AXI_read_addr = addr;
            temp_static_AXI_read_id = id;
            data_words_DIMS0 = data_words.size();
            temp_static_AXI_read_data_words = data_words;
            resp_DIMS0 = resp.size();
            temp_static_AXI_read_resp = resp;
            data_user_DIMS0 = data_user.size();
            temp_static_AXI_read_data_user = data_user;
            data_start_time_DIMS0 = data_start_time.size();
            temp_static_AXI_read_data_start_time = data_start_time;
            data_end_time_DIMS0 = data_end_time.size();
            temp_static_AXI_read_data_end_time = data_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            // In addition gets back updated sizes of unsized params.
            axi_AXI_read_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, data_words_DIMS0, resp_DIMS0, addr_user, data_user_DIMS0, address_to_data_latency, addr_start_time, addr_end_time, data_start_time_DIMS0, data_end_time_DIMS0, address_valid_delay, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_words.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_AXI_read_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_user.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, addr_user, address_to_data_latency, addr_start_time, addr_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_AXI_read_addr;
            id = temp_static_AXI_read_id;
            data_words = temp_static_AXI_read_data_words;
            temp_static_AXI_read_data_words.delete();
            resp = temp_static_AXI_read_resp;
            temp_static_AXI_read_resp.delete();
            data_user = temp_static_AXI_read_data_user;
            temp_static_AXI_read_data_user.delete();
            data_start_time = temp_static_AXI_read_data_start_time;
            temp_static_AXI_read_data_start_time.delete();
            data_end_time = temp_static_AXI_read_data_end_time;
            temp_static_AXI_read_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_AXI_read
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output int address_to_data_latency,
        output longint addr_start_time,
        output longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        output int address_valid_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_AXI_read_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, resp_DIMS0, data_user_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_words.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_AXI_read_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_user.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, addr_user, address_to_data_latency, addr_start_time, addr_end_time, address_valid_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_AXI_read_addr;
            id = temp_static_AXI_read_id;
            data_words = temp_static_AXI_read_data_words;
            temp_static_AXI_read_data_words.delete();
            resp = temp_static_AXI_read_resp;
            temp_static_AXI_read_resp.delete();
            data_user = temp_static_AXI_read_data_user;
            temp_static_AXI_read_data_user.delete();
            data_start_time = temp_static_AXI_read_data_start_time;
            temp_static_AXI_read_data_start_time.delete();
            data_end_time = temp_static_AXI_read_data_end_time;
            temp_static_AXI_read_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_AXI_write
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp,
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref int address_to_data_latency,
        ref int data_to_response_latency,
        ref int write_address_to_data_delay,
        ref int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        ref longint addr_start_time,
        ref longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        ref longint wr_resp_start_time,
        ref longint wr_resp_end_time,
        ref int address_valid_delay,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_AXI_write_addr = addr;
            temp_static_AXI_write_id = id;
            data_words_DIMS0 = data_words.size();
            temp_static_AXI_write_data_words = data_words;
            write_strobes_DIMS0 = write_strobes.size();
            temp_static_AXI_write_write_strobes = write_strobes;
            data_user_DIMS0 = data_user.size();
            temp_static_AXI_write_data_user = data_user;
            write_data_beats_delay_DIMS0 = write_data_beats_delay.size();
            temp_static_AXI_write_write_data_beats_delay = write_data_beats_delay;
            data_start_time_DIMS0 = data_start_time.size();
            temp_static_AXI_write_data_start_time = data_start_time;
            data_end_time_DIMS0 = data_end_time.size();
            temp_static_AXI_write_data_end_time = data_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            // In addition gets back updated sizes of unsized params.
            axi_AXI_write_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, data_words_DIMS0, write_strobes_DIMS0, resp, addr_user, data_user_DIMS0, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay_DIMS0, addr_start_time, addr_end_time, data_start_time_DIMS0, data_end_time_DIMS0, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_AXI_write_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_AXI_write_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_write_data_beats_delay.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, resp, addr_user, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, addr_start_time, addr_end_time, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_AXI_write_addr;
            id = temp_static_AXI_write_id;
            data_words = temp_static_AXI_write_data_words;
            temp_static_AXI_write_data_words.delete();
            write_strobes = temp_static_AXI_write_write_strobes;
            temp_static_AXI_write_write_strobes.delete();
            data_user = temp_static_AXI_write_data_user;
            temp_static_AXI_write_data_user.delete();
            write_data_beats_delay = temp_static_AXI_write_write_data_beats_delay;
            temp_static_AXI_write_write_data_beats_delay.delete();
            data_start_time = temp_static_AXI_write_data_start_time;
            temp_static_AXI_write_data_start_time.delete();
            data_end_time = temp_static_AXI_write_data_end_time;
            temp_static_AXI_write_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_AXI_write
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output axi_response_e resp,
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        output longint addr_start_time,
        output longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        output longint wr_resp_start_time,
        output longint wr_resp_end_time,
        output int address_valid_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_AXI_write_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_AXI_write_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_AXI_write_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_write_data_beats_delay.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, resp, addr_user, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, addr_start_time, addr_end_time, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_AXI_write_addr;
            id = temp_static_AXI_write_id;
            data_words = temp_static_AXI_write_data_words;
            temp_static_AXI_write_data_words.delete();
            write_strobes = temp_static_AXI_write_write_strobes;
            temp_static_AXI_write_write_strobes.delete();
            data_user = temp_static_AXI_write_data_user;
            temp_static_AXI_write_data_user.delete();
            write_data_beats_delay = temp_static_AXI_write_write_data_beats_delay;
            temp_static_AXI_write_write_data_beats_delay.delete();
            data_start_time = temp_static_AXI_write_data_start_time;
            temp_static_AXI_write_data_start_time.delete();
            data_end_time = temp_static_AXI_write_data_end_time;
            temp_static_AXI_write_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_data_resp
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref axi_response_e resp,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref longint data_start,
        ref longint data_end,
        ref longint response_start,
        ref int write_data_beats_delay[],
        ref longint data_beat_start_time[],
        ref longint data_beat_end_time[],
        ref longint response_end_time,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_beat_start_time_DIMS0;
                automatic int data_beat_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            data_words_DIMS0 = data_words.size();
            temp_static_data_resp_data_words = data_words;
            write_strobes_DIMS0 = write_strobes.size();
            temp_static_data_resp_write_strobes = write_strobes;
            temp_static_data_resp_id = id;
            data_user_DIMS0 = data_user.size();
            temp_static_data_resp_data_user = data_user;
            write_data_beats_delay_DIMS0 = write_data_beats_delay.size();
            temp_static_data_resp_write_data_beats_delay = write_data_beats_delay;
            data_beat_start_time_DIMS0 = data_beat_start_time.size();
            temp_static_data_resp_data_beat_start_time = data_beat_start_time;
            data_beat_end_time_DIMS0 = data_beat_end_time.size();
            temp_static_data_resp_data_beat_end_time = data_beat_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            // In addition gets back updated sizes of unsized params.
            axi_data_resp_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, data_words_DIMS0, write_strobes_DIMS0, resp, data_user_DIMS0, resp_user, data_start, data_end, response_start, write_data_beats_delay_DIMS0, data_beat_start_time_DIMS0, data_beat_end_time_DIMS0, response_end_time, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_data_resp_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_data_resp_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_data_resp_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_data_resp_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_data_resp_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_data_resp_write_data_beats_delay.delete();
            end
            if (data_beat_start_time_DIMS0 != 0)
            begin
                temp_static_data_resp_data_beat_start_time = new [data_beat_start_time_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_beat_start_time.delete();
            end
            if (data_beat_end_time_DIMS0 != 0)
            begin
                temp_static_data_resp_data_beat_end_time = new [data_beat_end_time_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_beat_end_time.delete();
            end
            // Call function to get the sized params
            axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, resp, resp_user, data_start, data_end, response_start, response_end_time, _unit_id); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data_words = temp_static_data_resp_data_words;
            temp_static_data_resp_data_words.delete();
            write_strobes = temp_static_data_resp_write_strobes;
            temp_static_data_resp_write_strobes.delete();
            id = temp_static_data_resp_id;
            data_user = temp_static_data_resp_data_user;
            temp_static_data_resp_data_user.delete();
            write_data_beats_delay = temp_static_data_resp_write_data_beats_delay;
            temp_static_data_resp_write_data_beats_delay.delete();
            data_beat_start_time = temp_static_data_resp_data_beat_start_time;
            temp_static_data_resp_data_beat_start_time.delete();
            data_beat_end_time = temp_static_data_resp_data_beat_end_time;
            temp_static_data_resp_data_beat_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_data_resp
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_response_e resp,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output longint data_start,
        output longint data_end,
        output longint response_start,
        ref int write_data_beats_delay[],
        ref longint data_beat_start_time[],
        ref longint data_beat_end_time[],
        output longint response_end_time,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_beat_start_time_DIMS0;
                automatic int data_beat_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_data_resp_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_beat_start_time_DIMS0, data_beat_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_data_resp_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_data_resp_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_data_resp_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_data_resp_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_data_resp_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_data_resp_write_data_beats_delay.delete();
            end
            if (data_beat_start_time_DIMS0 != 0)
            begin
                temp_static_data_resp_data_beat_start_time = new [data_beat_start_time_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_beat_start_time.delete();
            end
            if (data_beat_end_time_DIMS0 != 0)
            begin
                temp_static_data_resp_data_beat_end_time = new [data_beat_end_time_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_beat_end_time.delete();
            end
            // Call function to get the sized params
            axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, resp, resp_user, data_start, data_end, response_start, response_end_time, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data_words = temp_static_data_resp_data_words;
            temp_static_data_resp_data_words.delete();
            write_strobes = temp_static_data_resp_write_strobes;
            temp_static_data_resp_write_strobes.delete();
            id = temp_static_data_resp_id;
            data_user = temp_static_data_resp_data_user;
            temp_static_data_resp_data_user.delete();
            write_data_beats_delay = temp_static_data_resp_write_data_beats_delay;
            temp_static_data_resp_write_data_beats_delay.delete();
            data_beat_start_time = temp_static_data_resp_data_beat_start_time;
            temp_static_data_resp_data_beat_start_time.delete();
            data_beat_end_time = temp_static_data_resp_data_beat_end_time;
            temp_static_data_resp_data_beat_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            data_words_DIMS0 = data_words.size();
            temp_static_read_data_burst_data_words = data_words;
            resp_DIMS0 = resp.size();
            temp_static_read_data_burst_resp = resp;
            temp_static_read_data_burst_id = id;
            data_user_DIMS0 = data_user.size();
            temp_static_read_data_burst_data_user = data_user;
            data_start_time_DIMS0 = data_start_time.size();
            temp_static_read_data_burst_data_start_time = data_start_time;
            data_end_time_DIMS0 = data_end_time.size();
            temp_static_read_data_burst_data_end_time = data_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_data_burst_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, data_words_DIMS0, resp_DIMS0, data_user_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            temp_static_read_data_burst_data_words.delete();
            temp_static_read_data_burst_resp.delete();
            temp_static_read_data_burst_data_user.delete();
            temp_static_read_data_burst_data_start_time.delete();
            temp_static_read_data_burst_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, resp_DIMS0, data_user_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_read_data_burst_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_data_words.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_read_data_burst_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_read_data_burst_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_data_user.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_read_data_burst_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_read_data_burst_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data_words = temp_static_read_data_burst_data_words;
            temp_static_read_data_burst_data_words.delete();
            resp = temp_static_read_data_burst_resp;
            temp_static_read_data_burst_resp.delete();
            id = temp_static_read_data_burst_id;
            data_user = temp_static_read_data_burst_data_user;
            temp_static_read_data_burst_data_user.delete();
            data_start_time = temp_static_read_data_burst_data_start_time;
            temp_static_read_data_burst_data_start_time.delete();
            data_end_time = temp_static_read_data_burst_data_end_time;
            temp_static_read_data_burst_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref int write_data_beats_delay[],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            data_words_DIMS0 = data_words.size();
            temp_static_write_data_burst_data_words = data_words;
            write_strobes_DIMS0 = write_strobes.size();
            temp_static_write_data_burst_write_strobes = write_strobes;
            temp_static_write_data_burst_id = id;
            data_user_DIMS0 = data_user.size();
            temp_static_write_data_burst_data_user = data_user;
            write_data_beats_delay_DIMS0 = write_data_beats_delay.size();
            temp_static_write_data_burst_write_data_beats_delay = write_data_beats_delay;
            data_start_time_DIMS0 = data_start_time.size();
            temp_static_write_data_burst_data_start_time = data_start_time;
            data_end_time_DIMS0 = data_end_time.size();
            temp_static_write_data_burst_data_end_time = data_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_data_burst_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            temp_static_write_data_burst_data_words.delete();
            temp_static_write_data_burst_write_strobes.delete();
            temp_static_write_data_burst_data_user.delete();
            temp_static_write_data_burst_write_data_beats_delay.delete();
            temp_static_write_data_burst_data_start_time.delete();
            temp_static_write_data_burst_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref int write_data_beats_delay[],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_write_data_burst_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_write_data_burst_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_write_data_burst_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_write_data_burst_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_write_data_beats_delay.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_write_data_burst_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_write_data_burst_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data_words = temp_static_write_data_burst_data_words;
            temp_static_write_data_burst_data_words.delete();
            write_strobes = temp_static_write_data_burst_write_strobes;
            temp_static_write_data_burst_write_strobes.delete();
            id = temp_static_write_data_burst_id;
            data_user = temp_static_write_data_burst_data_user;
            temp_static_write_data_burst_data_user.delete();
            write_data_beats_delay = temp_static_write_data_burst_write_data_beats_delay;
            temp_static_write_data_burst_write_data_beats_delay.delete();
            data_start_time = temp_static_write_data_burst_data_start_time;
            temp_static_write_data_burst_data_start_time.delete();
            data_end_time = temp_static_write_data_burst_data_end_time;
            temp_static_write_data_burst_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_read_addr_channel_phase_addr = addr;
            temp_static_read_addr_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_addr_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, size, burst, lock, cache, prot, addr_user, address_valid_delay, address_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_read_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, size, burst, lock, cache, prot, addr_user, address_valid_delay, address_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_read_addr_channel_phase_addr;
            id = temp_static_read_addr_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_read_channel_phase_data = data;
            temp_static_read_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, resp, data_user, data_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_read_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, last, resp, data_user, data_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data = temp_static_read_channel_phase_data;
            id = temp_static_read_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_addr_channel_phase_addr = addr;
            temp_static_write_addr_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_addr_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, size, burst, lock, cache, prot, addr_user, address_valid_delay, address_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, size, burst, lock, cache, prot, addr_user, address_valid_delay, address_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_write_addr_channel_phase_addr;
            id = temp_static_write_addr_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_channel_phase_data = data;
            temp_static_write_channel_phase_write_strobes = write_strobes;
            temp_static_write_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, data_user, data_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, last, data_user, data_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data = temp_static_write_channel_phase_data;
            write_strobes = temp_static_write_channel_phase_write_strobes;
            id = temp_static_write_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_resp_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int write_response_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_resp_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_resp_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, resp, resp_user, write_response_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_resp_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        output int write_response_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_resp_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, resp, resp_user, write_response_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            id = temp_static_write_resp_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_read_addr_channel_cycle_addr = addr;
            temp_static_read_addr_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, size, burst, lock, cache, prot, addr_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_read_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, size, burst, lock, cache, prot, addr_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_read_addr_channel_cycle_addr;
            id = temp_static_read_addr_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_read_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_read_channel_cycle_data = data;
            temp_static_read_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, resp, data_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_read_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, last, resp, data_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data = temp_static_read_channel_cycle_data;
            id = temp_static_read_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_addr_channel_cycle_addr = addr;
            temp_static_write_addr_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, size, burst, lock, cache, prot, addr_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, size, burst, lock, cache, prot, addr_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_write_addr_channel_cycle_addr;
            id = temp_static_write_addr_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_channel_cycle_data = data;
            temp_static_write_channel_cycle_strb = strb;
            temp_static_write_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, data_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, last, data_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data = temp_static_write_channel_cycle_data;
            strb = temp_static_write_channel_cycle_strb;
            id = temp_static_write_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_resp_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_resp_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, resp, resp_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_resp_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_resp_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, resp, resp_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            id = temp_static_write_resp_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_resp_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_resp_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask


    //-------------------------------------------------------------------------
    // Generic Interface Configuration Support
    //

    import "DPI-C" context axi_set_interface = function void axi_set_interface
    (
        input int what,
        input int arg1,
        input int arg2,
        input int arg3,
        input int arg4,
        input int arg5,
        input int arg6,
        input int arg7,
        input int arg8,
        input int arg9,
        input int arg10
    );
    import "DPI-C" context axi_get_interface = function int axi_get_interface
    (
        input int what,
        input int arg1,
        input int arg2,
        input int arg3,
        input int arg4,
        input int arg5,
        input int arg6,
        input int arg7,
        input int arg8,
        input int arg9
    );


    //-------------------------------------------------------------------------
    // Functions to get the hierarchic name of this interface
    //
    import "DPI-C" context axi_get_full_name = function string axi_get_full_name();


    //-------------------------------------------------------------------------
    // Abstraction level Support
    //

    import "DPI-C" context axi_set_master_end_abstraction_level =
    function void axi_set_master_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_master_end_abstraction_level =
    function void axi_get_master_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_slave_end_abstraction_level =
    function void axi_set_slave_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_slave_end_abstraction_level =
    function void axi_get_slave_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_clock_source_end_abstraction_level =
    function void axi_set_clock_source_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_clock_source_end_abstraction_level =
    function void axi_get_clock_source_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_reset_source_end_abstraction_level =
    function void axi_set_reset_source_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_reset_source_end_abstraction_level =
    function void axi_get_reset_source_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );

    //-------------------------------------------------------------------------
    // Wire Level Interface Support
    //
    logic internal_ACLK = 'z;
    logic internal_ARESETn = 'z;
    logic internal_AWVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  internal_AWADDR = 'z;
    logic [3:0] internal_AWLEN = 'z;
    logic [2:0] internal_AWSIZE = 'z;
    logic [1:0] internal_AWBURST = 'z;
    logic [1:0] internal_AWLOCK = 'z;
    logic [3:0] internal_AWCACHE = 'z;
    logic [2:0] internal_AWPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_AWID = 'z;
    logic internal_AWREADY = 'z;
    logic [7:0] internal_AWUSER = 'z;
    logic internal_ARVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  internal_ARADDR = 'z;
    logic [3:0] internal_ARLEN = 'z;
    logic [2:0] internal_ARSIZE = 'z;
    logic [1:0] internal_ARBURST = 'z;
    logic [1:0] internal_ARLOCK = 'z;
    logic [3:0] internal_ARCACHE = 'z;
    logic [2:0] internal_ARPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_ARID = 'z;
    logic internal_ARREADY = 'z;
    logic [7:0] internal_ARUSER = 'z;
    logic internal_RVALID = 'z;
    logic internal_RLAST = 'z;
    logic [((AXI_RDATA_WIDTH) - 1):0]  internal_RDATA = 'z;
    logic [1:0] internal_RRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_RID = 'z;
    logic internal_RREADY = 'z;
    logic [7:0] internal_RUSER = 'z;
    logic internal_WVALID = 'z;
    logic internal_WLAST = 'z;
    logic [((AXI_WDATA_WIDTH) - 1):0]  internal_WDATA = 'z;
    logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  internal_WSTRB = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_WID = 'z;
    logic internal_WREADY = 'z;
    logic [7:0] internal_WUSER = 'z;
    logic internal_BVALID = 'z;
    logic [1:0] internal_BRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_BID = 'z;
    logic internal_BREADY = 'z;
    logic [7:0] internal_BUSER = 'z;

    import "DPI-C" context function void axi_set_ACLK_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit ACLK_param
    );
    import "DPI-C" context function void axi_propagate_ACLK_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ACLK_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit ACLK_param

    );
    export "DPI-C" function axi_initialise_ACLK_from_CY;

    import "DPI-C" context function void axi_set_ARESETn_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARESETn_param
    );
    import "DPI-C" context function void axi_propagate_ARESETn_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARESETn_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARESETn_param

    );
    export "DPI-C" function axi_initialise_ARESETn_from_CY;

    import "DPI-C" context function void axi_set_AWVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic AWVALID_param
    );
    import "DPI-C" context function void axi_propagate_AWVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic AWVALID_param

    );
    export "DPI-C" function axi_initialise_AWVALID_from_CY;

    import "DPI-C" context function void axi_set_AWADDR_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  AWADDR_param
    );
    import "DPI-C" context function void axi_propagate_AWADDR_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWADDR_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_AWADDR_from_CY_index1;
    export "DPI-C" function axi_initialise_AWADDR_from_CY;

    import "DPI-C" context function void axi_set_AWLEN_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] AWLEN_param
    );
    import "DPI-C" context function void axi_propagate_AWLEN_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWLEN_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] AWLEN_param

    );
    export "DPI-C" function axi_initialise_AWLEN_from_CY;

    import "DPI-C" context function void axi_set_AWSIZE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] AWSIZE_param
    );
    import "DPI-C" context function void axi_propagate_AWSIZE_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWSIZE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] AWSIZE_param

    );
    export "DPI-C" function axi_initialise_AWSIZE_from_CY;

    import "DPI-C" context function void axi_set_AWBURST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] AWBURST_param
    );
    import "DPI-C" context function void axi_propagate_AWBURST_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWBURST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] AWBURST_param

    );
    export "DPI-C" function axi_initialise_AWBURST_from_CY;

    import "DPI-C" context function void axi_set_AWLOCK_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] AWLOCK_param
    );
    import "DPI-C" context function void axi_propagate_AWLOCK_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWLOCK_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] AWLOCK_param

    );
    export "DPI-C" function axi_initialise_AWLOCK_from_CY;

    import "DPI-C" context function void axi_set_AWCACHE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] AWCACHE_param
    );
    import "DPI-C" context function void axi_propagate_AWCACHE_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWCACHE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] AWCACHE_param

    );
    export "DPI-C" function axi_initialise_AWCACHE_from_CY;

    import "DPI-C" context function void axi_set_AWPROT_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] AWPROT_param
    );
    import "DPI-C" context function void axi_propagate_AWPROT_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWPROT_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] AWPROT_param

    );
    export "DPI-C" function axi_initialise_AWPROT_from_CY;

    import "DPI-C" context function void axi_set_AWID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  AWID_param
    );
    import "DPI-C" context function void axi_propagate_AWID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_AWID_from_CY_index1;
    export "DPI-C" function axi_initialise_AWID_from_CY;

    import "DPI-C" context function void axi_set_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic AWREADY_param
    );
    import "DPI-C" context function void axi_propagate_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic AWREADY_param

    );
    export "DPI-C" function axi_initialise_AWREADY_from_CY;

    import "DPI-C" context function void axi_set_AWUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] AWUSER_param
    );
    import "DPI-C" context function void axi_propagate_AWUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] AWUSER_param

    );
    export "DPI-C" function axi_initialise_AWUSER_from_CY;

    import "DPI-C" context function void axi_set_ARVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARVALID_param
    );
    import "DPI-C" context function void axi_propagate_ARVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARVALID_param

    );
    export "DPI-C" function axi_initialise_ARVALID_from_CY;

    import "DPI-C" context function void axi_set_ARADDR_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  ARADDR_param
    );
    import "DPI-C" context function void axi_propagate_ARADDR_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARADDR_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_ARADDR_from_CY_index1;
    export "DPI-C" function axi_initialise_ARADDR_from_CY;

    import "DPI-C" context function void axi_set_ARLEN_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] ARLEN_param
    );
    import "DPI-C" context function void axi_propagate_ARLEN_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARLEN_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] ARLEN_param

    );
    export "DPI-C" function axi_initialise_ARLEN_from_CY;

    import "DPI-C" context function void axi_set_ARSIZE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] ARSIZE_param
    );
    import "DPI-C" context function void axi_propagate_ARSIZE_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARSIZE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] ARSIZE_param

    );
    export "DPI-C" function axi_initialise_ARSIZE_from_CY;

    import "DPI-C" context function void axi_set_ARBURST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] ARBURST_param
    );
    import "DPI-C" context function void axi_propagate_ARBURST_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARBURST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] ARBURST_param

    );
    export "DPI-C" function axi_initialise_ARBURST_from_CY;

    import "DPI-C" context function void axi_set_ARLOCK_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] ARLOCK_param
    );
    import "DPI-C" context function void axi_propagate_ARLOCK_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARLOCK_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] ARLOCK_param

    );
    export "DPI-C" function axi_initialise_ARLOCK_from_CY;

    import "DPI-C" context function void axi_set_ARCACHE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] ARCACHE_param
    );
    import "DPI-C" context function void axi_propagate_ARCACHE_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARCACHE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] ARCACHE_param

    );
    export "DPI-C" function axi_initialise_ARCACHE_from_CY;

    import "DPI-C" context function void axi_set_ARPROT_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] ARPROT_param
    );
    import "DPI-C" context function void axi_propagate_ARPROT_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARPROT_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] ARPROT_param

    );
    export "DPI-C" function axi_initialise_ARPROT_from_CY;

    import "DPI-C" context function void axi_set_ARID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  ARID_param
    );
    import "DPI-C" context function void axi_propagate_ARID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_ARID_from_CY_index1;
    export "DPI-C" function axi_initialise_ARID_from_CY;

    import "DPI-C" context function void axi_set_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARREADY_param
    );
    import "DPI-C" context function void axi_propagate_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARREADY_param

    );
    export "DPI-C" function axi_initialise_ARREADY_from_CY;

    import "DPI-C" context function void axi_set_ARUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] ARUSER_param
    );
    import "DPI-C" context function void axi_propagate_ARUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] ARUSER_param

    );
    export "DPI-C" function axi_initialise_ARUSER_from_CY;

    import "DPI-C" context function void axi_set_RVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RVALID_param
    );
    import "DPI-C" context function void axi_propagate_RVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RVALID_param

    );
    export "DPI-C" function axi_initialise_RVALID_from_CY;

    import "DPI-C" context function void axi_set_RLAST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RLAST_param
    );
    import "DPI-C" context function void axi_propagate_RLAST_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RLAST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RLAST_param

    );
    export "DPI-C" function axi_initialise_RLAST_from_CY;

    import "DPI-C" context function void axi_set_RDATA_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  RDATA_param
    );
    import "DPI-C" context function void axi_propagate_RDATA_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RDATA_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_RDATA_from_CY_index1;
    export "DPI-C" function axi_initialise_RDATA_from_CY;

    import "DPI-C" context function void axi_set_RRESP_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] RRESP_param
    );
    import "DPI-C" context function void axi_propagate_RRESP_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RRESP_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] RRESP_param

    );
    export "DPI-C" function axi_initialise_RRESP_from_CY;

    import "DPI-C" context function void axi_set_RID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  RID_param
    );
    import "DPI-C" context function void axi_propagate_RID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_RID_from_CY_index1;
    export "DPI-C" function axi_initialise_RID_from_CY;

    import "DPI-C" context function void axi_set_RREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RREADY_param
    );
    import "DPI-C" context function void axi_propagate_RREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RREADY_param

    );
    export "DPI-C" function axi_initialise_RREADY_from_CY;

    import "DPI-C" context function void axi_set_RUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] RUSER_param
    );
    import "DPI-C" context function void axi_propagate_RUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] RUSER_param

    );
    export "DPI-C" function axi_initialise_RUSER_from_CY;

    import "DPI-C" context function void axi_set_WVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WVALID_param
    );
    import "DPI-C" context function void axi_propagate_WVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WVALID_param

    );
    export "DPI-C" function axi_initialise_WVALID_from_CY;

    import "DPI-C" context function void axi_set_WLAST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WLAST_param
    );
    import "DPI-C" context function void axi_propagate_WLAST_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WLAST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WLAST_param

    );
    export "DPI-C" function axi_initialise_WLAST_from_CY;

    import "DPI-C" context function void axi_set_WDATA_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  WDATA_param
    );
    import "DPI-C" context function void axi_propagate_WDATA_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WDATA_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_WDATA_from_CY_index1;
    export "DPI-C" function axi_initialise_WDATA_from_CY;

    import "DPI-C" context function void axi_set_WSTRB_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  WSTRB_param
    );
    import "DPI-C" context function void axi_propagate_WSTRB_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WSTRB_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_WSTRB_from_CY_index1;
    export "DPI-C" function axi_initialise_WSTRB_from_CY;

    import "DPI-C" context function void axi_set_WID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  WID_param
    );
    import "DPI-C" context function void axi_propagate_WID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_WID_from_CY_index1;
    export "DPI-C" function axi_initialise_WID_from_CY;

    import "DPI-C" context function void axi_set_WREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WREADY_param
    );
    import "DPI-C" context function void axi_propagate_WREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WREADY_param

    );
    export "DPI-C" function axi_initialise_WREADY_from_CY;

    import "DPI-C" context function void axi_set_WUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] WUSER_param
    );
    import "DPI-C" context function void axi_propagate_WUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] WUSER_param

    );
    export "DPI-C" function axi_initialise_WUSER_from_CY;

    import "DPI-C" context function void axi_set_BVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic BVALID_param
    );
    import "DPI-C" context function void axi_propagate_BVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic BVALID_param

    );
    export "DPI-C" function axi_initialise_BVALID_from_CY;

    import "DPI-C" context function void axi_set_BRESP_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] BRESP_param
    );
    import "DPI-C" context function void axi_propagate_BRESP_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BRESP_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] BRESP_param

    );
    export "DPI-C" function axi_initialise_BRESP_from_CY;

    import "DPI-C" context function void axi_set_BID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  BID_param
    );
    import "DPI-C" context function void axi_propagate_BID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_BID_from_CY_index1;
    export "DPI-C" function axi_initialise_BID_from_CY;

    import "DPI-C" context function void axi_set_BREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic BREADY_param
    );
    import "DPI-C" context function void axi_propagate_BREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic BREADY_param

    );
    export "DPI-C" function axi_initialise_BREADY_from_CY;

    import "DPI-C" context function void axi_set_BUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] BUSER_param
    );
    import "DPI-C" context function void axi_propagate_BUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] BUSER_param

    );
    export "DPI-C" function axi_initialise_BUSER_from_CY;

    import "DPI-C" context function void axi_set_config_write_ctrl_to_data_mintime_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_write_ctrl_to_data_mintime_param
    );
    import "DPI-C" context function void axi_propagate_config_write_ctrl_to_data_mintime_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_write_ctrl_to_data_mintime_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_write_ctrl_to_data_mintime_param

    );
    export "DPI-C" function axi_set_config_write_ctrl_to_data_mintime_from_CY;

    import "DPI-C" context function void axi_set_config_master_write_delay_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_master_write_delay_param
    );
    import "DPI-C" context function void axi_propagate_config_master_write_delay_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_deprecated_config_master_write_delay_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_master_write_delay_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_master_write_delay_param

    );
    export "DPI-C" function axi_set_config_master_write_delay_from_CY;

    import "DPI-C" context function void axi_set_config_enable_all_assertions_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_enable_all_assertions_param
    );
    import "DPI-C" context function void axi_propagate_config_enable_all_assertions_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_enable_all_assertions_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_enable_all_assertions_param

    );
    export "DPI-C" function axi_set_config_enable_all_assertions_from_CY;

    import "DPI-C" context function void axi_set_config_enable_assertion_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param
    );
    import "DPI-C" context function void axi_propagate_config_enable_assertion_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_enable_assertion_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param

    );
    export "DPI-C" function axi_set_config_enable_assertion_from_CY;

    import "DPI-C" context function void axi_set_config_slave_start_addr_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input bit  config_slave_start_addr_param
    );
    import "DPI-C" context function void axi_propagate_config_slave_start_addr_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_deprecated_config_slave_start_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_slave_start_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_config_slave_start_addr_from_CY_index1;

    import "DPI-C" context function void axi_set_config_slave_end_addr_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input bit  config_slave_end_addr_param
    );
    import "DPI-C" context function void axi_propagate_config_slave_end_addr_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_deprecated_config_slave_end_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_slave_end_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_config_slave_end_addr_from_CY_index1;

    import "DPI-C" context function void axi_set_config_support_exclusive_access_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_support_exclusive_access_param
    );
    import "DPI-C" context function void axi_propagate_config_support_exclusive_access_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_support_exclusive_access_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_support_exclusive_access_param

    );
    export "DPI-C" function axi_set_config_support_exclusive_access_from_CY;

    import "DPI-C" context function void axi_set_config_read_data_reordering_depth_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_read_data_reordering_depth_param
    );
    import "DPI-C" context function void axi_propagate_config_read_data_reordering_depth_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_read_data_reordering_depth_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_read_data_reordering_depth_param

    );
    export "DPI-C" function axi_set_config_read_data_reordering_depth_from_CY;

    import "DPI-C" context function void axi_set_config_max_transaction_time_factor_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_transaction_time_factor_param
    );
    import "DPI-C" context function void axi_propagate_config_max_transaction_time_factor_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_transaction_time_factor_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_transaction_time_factor_param

    );
    export "DPI-C" function axi_set_config_max_transaction_time_factor_from_CY;

    import "DPI-C" context function void axi_set_config_timeout_max_data_transfer_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_timeout_max_data_transfer_param
    );
    import "DPI-C" context function void axi_propagate_config_timeout_max_data_transfer_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_timeout_max_data_transfer_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_timeout_max_data_transfer_param

    );
    export "DPI-C" function axi_set_config_timeout_max_data_transfer_from_CY;

    import "DPI-C" context function void axi_set_config_burst_timeout_factor_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_burst_timeout_factor_param
    );
    import "DPI-C" context function void axi_propagate_config_burst_timeout_factor_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_burst_timeout_factor_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_burst_timeout_factor_param

    );
    export "DPI-C" function axi_set_config_burst_timeout_factor_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_AWVALID_assertion_to_AWREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_ARVALID_assertion_to_ARREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_RVALID_assertion_to_RREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_RVALID_assertion_to_RREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_RVALID_assertion_to_RREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_BVALID_assertion_to_BREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_BVALID_assertion_to_BREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_BVALID_assertion_to_BREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_WVALID_assertion_to_WREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_WVALID_assertion_to_WREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_WVALID_assertion_to_WREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_CY;

    import "DPI-C" context function void axi_set_config_master_error_position_from_SystemVerilog
    (
        input longint _iface_ref,
        input axi_error_e config_master_error_position_param
    );
    import "DPI-C" context function void axi_propagate_config_master_error_position_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_deprecated_config_master_error_position_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_master_error_position_into_SystemVerilog
    (
        input longint _iface_ref,
        output axi_error_e config_master_error_position_param

    );
    export "DPI-C" function axi_set_config_master_error_position_from_CY;

    import "DPI-C" context function void axi_set_config_setup_time_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_setup_time_param
    );
    import "DPI-C" context function void axi_propagate_config_setup_time_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_setup_time_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_setup_time_param

    );
    export "DPI-C" function axi_set_config_setup_time_from_CY;

    import "DPI-C" context function void axi_set_config_hold_time_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_hold_time_param
    );
    import "DPI-C" context function void axi_propagate_config_hold_time_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_hold_time_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_hold_time_param

    );
    export "DPI-C" function axi_set_config_hold_time_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_wr_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_wr_param
    );
    import "DPI-C" context function void axi_propagate_config_max_outstanding_wr_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_outstanding_wr_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_wr_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_wr_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_rd_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_rd_param
    );
    import "DPI-C" context function void axi_propagate_config_max_outstanding_rd_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_outstanding_rd_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_rd_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_rd_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_rw_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_rw_param
    );
    import "DPI-C" context function void axi_propagate_config_max_outstanding_rw_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_outstanding_rw_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_rw_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_rw_from_CY;

    import "DPI-C" context function void axi_set_config_is_issuing_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_is_issuing_param
    );
    import "DPI-C" context function void axi_propagate_config_is_issuing_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_is_issuing_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_is_issuing_param

    );
    export "DPI-C" function axi_set_config_is_issuing_from_CY;

    function void axi_initialise_ACLK_from_CY();
        internal_ACLK = 'z;
        m_ACLK = 'z;
    endfunction

    function void axi_initialise_ARESETn_from_CY();
        internal_ARESETn = 'z;
        m_ARESETn = 'z;
    endfunction

    function void axi_initialise_AWVALID_from_CY();
        internal_AWVALID = 'z;
        m_AWVALID = 'z;
    endfunction

    function void axi_set_AWADDR_from_CY_index1( int _this_dot_1, logic  AWADDR_param );
        internal_AWADDR[_this_dot_1] = AWADDR_param;
    endfunction

    function void axi_initialise_AWADDR_from_CY();
        internal_AWADDR = 'z;
        m_AWADDR = 'z;
    endfunction

    function void axi_initialise_AWLEN_from_CY();
        internal_AWLEN = 'z;
        m_AWLEN = 'z;
    endfunction

    function void axi_initialise_AWSIZE_from_CY();
        internal_AWSIZE = 'z;
        m_AWSIZE = 'z;
    endfunction

    function void axi_initialise_AWBURST_from_CY();
        internal_AWBURST = 'z;
        m_AWBURST = 'z;
    endfunction

    function void axi_initialise_AWLOCK_from_CY();
        internal_AWLOCK = 'z;
        m_AWLOCK = 'z;
    endfunction

    function void axi_initialise_AWCACHE_from_CY();
        internal_AWCACHE = 'z;
        m_AWCACHE = 'z;
    endfunction

    function void axi_initialise_AWPROT_from_CY();
        internal_AWPROT = 'z;
        m_AWPROT = 'z;
    endfunction

    function void axi_set_AWID_from_CY_index1( int _this_dot_1, logic  AWID_param );
        internal_AWID[_this_dot_1] = AWID_param;
    endfunction

    function void axi_initialise_AWID_from_CY();
        internal_AWID = 'z;
        m_AWID = 'z;
    endfunction

    function void axi_initialise_AWREADY_from_CY();
        internal_AWREADY = 'z;
        m_AWREADY = 'z;
    endfunction

    function void axi_initialise_AWUSER_from_CY();
        internal_AWUSER = 'z;
        m_AWUSER = 'z;
    endfunction

    function void axi_initialise_ARVALID_from_CY();
        internal_ARVALID = 'z;
        m_ARVALID = 'z;
    endfunction

    function void axi_set_ARADDR_from_CY_index1( int _this_dot_1, logic  ARADDR_param );
        internal_ARADDR[_this_dot_1] = ARADDR_param;
    endfunction

    function void axi_initialise_ARADDR_from_CY();
        internal_ARADDR = 'z;
        m_ARADDR = 'z;
    endfunction

    function void axi_initialise_ARLEN_from_CY();
        internal_ARLEN = 'z;
        m_ARLEN = 'z;
    endfunction

    function void axi_initialise_ARSIZE_from_CY();
        internal_ARSIZE = 'z;
        m_ARSIZE = 'z;
    endfunction

    function void axi_initialise_ARBURST_from_CY();
        internal_ARBURST = 'z;
        m_ARBURST = 'z;
    endfunction

    function void axi_initialise_ARLOCK_from_CY();
        internal_ARLOCK = 'z;
        m_ARLOCK = 'z;
    endfunction

    function void axi_initialise_ARCACHE_from_CY();
        internal_ARCACHE = 'z;
        m_ARCACHE = 'z;
    endfunction

    function void axi_initialise_ARPROT_from_CY();
        internal_ARPROT = 'z;
        m_ARPROT = 'z;
    endfunction

    function void axi_set_ARID_from_CY_index1( int _this_dot_1, logic  ARID_param );
        internal_ARID[_this_dot_1] = ARID_param;
    endfunction

    function void axi_initialise_ARID_from_CY();
        internal_ARID = 'z;
        m_ARID = 'z;
    endfunction

    function void axi_initialise_ARREADY_from_CY();
        internal_ARREADY = 'z;
        m_ARREADY = 'z;
    endfunction

    function void axi_initialise_ARUSER_from_CY();
        internal_ARUSER = 'z;
        m_ARUSER = 'z;
    endfunction

    function void axi_initialise_RVALID_from_CY();
        internal_RVALID = 'z;
        m_RVALID = 'z;
    endfunction

    function void axi_initialise_RLAST_from_CY();
        internal_RLAST = 'z;
        m_RLAST = 'z;
    endfunction

    function void axi_set_RDATA_from_CY_index1( int _this_dot_1, logic  RDATA_param );
        internal_RDATA[_this_dot_1] = RDATA_param;
    endfunction

    function void axi_initialise_RDATA_from_CY();
        internal_RDATA = 'z;
        m_RDATA = 'z;
    endfunction

    function void axi_initialise_RRESP_from_CY();
        internal_RRESP = 'z;
        m_RRESP = 'z;
    endfunction

    function void axi_set_RID_from_CY_index1( int _this_dot_1, logic  RID_param );
        internal_RID[_this_dot_1] = RID_param;
    endfunction

    function void axi_initialise_RID_from_CY();
        internal_RID = 'z;
        m_RID = 'z;
    endfunction

    function void axi_initialise_RREADY_from_CY();
        internal_RREADY = 'z;
        m_RREADY = 'z;
    endfunction

    function void axi_initialise_RUSER_from_CY();
        internal_RUSER = 'z;
        m_RUSER = 'z;
    endfunction

    function void axi_initialise_WVALID_from_CY();
        internal_WVALID = 'z;
        m_WVALID = 'z;
    endfunction

    function void axi_initialise_WLAST_from_CY();
        internal_WLAST = 'z;
        m_WLAST = 'z;
    endfunction

    function void axi_set_WDATA_from_CY_index1( int _this_dot_1, logic  WDATA_param );
        internal_WDATA[_this_dot_1] = WDATA_param;
    endfunction

    function void axi_initialise_WDATA_from_CY();
        internal_WDATA = 'z;
        m_WDATA = 'z;
    endfunction

    function void axi_set_WSTRB_from_CY_index1( int _this_dot_1, logic  WSTRB_param );
        internal_WSTRB[_this_dot_1] = WSTRB_param;
    endfunction

    function void axi_initialise_WSTRB_from_CY();
        internal_WSTRB = 'z;
        m_WSTRB = 'z;
    endfunction

    function void axi_set_WID_from_CY_index1( int _this_dot_1, logic  WID_param );
        internal_WID[_this_dot_1] = WID_param;
    endfunction

    function void axi_initialise_WID_from_CY();
        internal_WID = 'z;
        m_WID = 'z;
    endfunction

    function void axi_initialise_WREADY_from_CY();
        internal_WREADY = 'z;
        m_WREADY = 'z;
    endfunction

    function void axi_initialise_WUSER_from_CY();
        internal_WUSER = 'z;
        m_WUSER = 'z;
    endfunction

    function void axi_initialise_BVALID_from_CY();
        internal_BVALID = 'z;
        m_BVALID = 'z;
    endfunction

    function void axi_initialise_BRESP_from_CY();
        internal_BRESP = 'z;
        m_BRESP = 'z;
    endfunction

    function void axi_set_BID_from_CY_index1( int _this_dot_1, logic  BID_param );
        internal_BID[_this_dot_1] = BID_param;
    endfunction

    function void axi_initialise_BID_from_CY();
        internal_BID = 'z;
        m_BID = 'z;
    endfunction

    function void axi_initialise_BREADY_from_CY();
        internal_BREADY = 'z;
        m_BREADY = 'z;
    endfunction

    function void axi_initialise_BUSER_from_CY();
        internal_BUSER = 'z;
        m_BUSER = 'z;
    endfunction

    function void axi_set_config_write_ctrl_to_data_mintime_from_CY( int unsigned config_write_ctrl_to_data_mintime_param );
        config_write_ctrl_to_data_mintime = config_write_ctrl_to_data_mintime_param;
    endfunction

    function void axi_set_config_master_write_delay_from_CY( bit config_master_write_delay_param );
        config_master_write_delay = config_master_write_delay_param;
    endfunction

    function void axi_set_config_enable_all_assertions_from_CY( bit config_enable_all_assertions_param );
        config_enable_all_assertions = config_enable_all_assertions_param;
    endfunction

    function void axi_set_config_enable_assertion_from_CY( bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
        config_enable_assertion = config_enable_assertion_param;
    endfunction

    function void axi_set_config_slave_start_addr_from_CY_index1( int _this_dot_1, bit  config_slave_start_addr_param );
        config_slave_start_addr[_this_dot_1] = config_slave_start_addr_param;
    endfunction

    function void axi_set_config_slave_end_addr_from_CY_index1( int _this_dot_1, bit  config_slave_end_addr_param );
        config_slave_end_addr[_this_dot_1] = config_slave_end_addr_param;
    endfunction

    function void axi_set_config_support_exclusive_access_from_CY( bit config_support_exclusive_access_param );
        config_support_exclusive_access = config_support_exclusive_access_param;
    endfunction

    function void axi_set_config_read_data_reordering_depth_from_CY( int unsigned config_read_data_reordering_depth_param );
        config_read_data_reordering_depth = config_read_data_reordering_depth_param;
    endfunction

    function void axi_set_config_max_transaction_time_factor_from_CY( int unsigned config_max_transaction_time_factor_param );
        config_max_transaction_time_factor = config_max_transaction_time_factor_param;
    endfunction

    function void axi_set_config_timeout_max_data_transfer_from_CY( int config_timeout_max_data_transfer_param );
        config_timeout_max_data_transfer = config_timeout_max_data_transfer_param;
    endfunction

    function void axi_set_config_burst_timeout_factor_from_CY( int unsigned config_burst_timeout_factor_param );
        config_burst_timeout_factor = config_burst_timeout_factor_param;
    endfunction

    function void axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_CY( int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
        config_max_latency_AWVALID_assertion_to_AWREADY = config_max_latency_AWVALID_assertion_to_AWREADY_param;
    endfunction

    function void axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_CY( int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
        config_max_latency_ARVALID_assertion_to_ARREADY = config_max_latency_ARVALID_assertion_to_ARREADY_param;
    endfunction

    function void axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_CY( int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
        config_max_latency_RVALID_assertion_to_RREADY = config_max_latency_RVALID_assertion_to_RREADY_param;
    endfunction

    function void axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_CY( int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
        config_max_latency_BVALID_assertion_to_BREADY = config_max_latency_BVALID_assertion_to_BREADY_param;
    endfunction

    function void axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_CY( int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
        config_max_latency_WVALID_assertion_to_WREADY = config_max_latency_WVALID_assertion_to_WREADY_param;
    endfunction

    function void axi_set_config_master_error_position_from_CY( axi_error_e config_master_error_position_param );
        config_master_error_position = config_master_error_position_param;
    endfunction

    function void axi_set_config_setup_time_from_CY( int config_setup_time_param );
        config_setup_time = config_setup_time_param;
    endfunction

    function void axi_set_config_hold_time_from_CY( int config_hold_time_param );
        config_hold_time = config_hold_time_param;
    endfunction

    function void axi_set_config_max_outstanding_wr_from_CY( int config_max_outstanding_wr_param );
        config_max_outstanding_wr = config_max_outstanding_wr_param;
    endfunction

    function void axi_set_config_max_outstanding_rd_from_CY( int config_max_outstanding_rd_param );
        config_max_outstanding_rd = config_max_outstanding_rd_param;
    endfunction

    function void axi_set_config_max_outstanding_rw_from_CY( int config_max_outstanding_rw_param );
        config_max_outstanding_rw = config_max_outstanding_rw_param;
    endfunction

    function void axi_set_config_is_issuing_from_CY( bit config_is_issuing_param );
        config_is_issuing = config_is_issuing_param;
    endfunction



    //--------------------------------------------------------------------------
    //
    // Group:- TLM Interface Support
    //
    //--------------------------------------------------------------------------
    export "DPI-C" axi_get_temp_static_rw_transaction_addr = function axi_get_temp_static_rw_transaction_addr;
    export "DPI-C" axi_set_temp_static_rw_transaction_addr = function axi_set_temp_static_rw_transaction_addr;
    export "DPI-C" axi_get_temp_static_rw_transaction_id = function axi_get_temp_static_rw_transaction_id;
    export "DPI-C" axi_set_temp_static_rw_transaction_id = function axi_set_temp_static_rw_transaction_id;
    export "DPI-C" axi_get_temp_static_rw_transaction_data_words = function axi_get_temp_static_rw_transaction_data_words;
    export "DPI-C" axi_set_temp_static_rw_transaction_data_words = function axi_set_temp_static_rw_transaction_data_words;
    export "DPI-C" axi_get_temp_static_rw_transaction_write_strobes = function axi_get_temp_static_rw_transaction_write_strobes;
    export "DPI-C" axi_set_temp_static_rw_transaction_write_strobes = function axi_set_temp_static_rw_transaction_write_strobes;
    export "DPI-C" axi_get_temp_static_rw_transaction_resp = function axi_get_temp_static_rw_transaction_resp;
    export "DPI-C" axi_set_temp_static_rw_transaction_resp = function axi_set_temp_static_rw_transaction_resp;
    export "DPI-C" axi_get_temp_static_rw_transaction_data_user = function axi_get_temp_static_rw_transaction_data_user;
    export "DPI-C" axi_set_temp_static_rw_transaction_data_user = function axi_set_temp_static_rw_transaction_data_user;
    export "DPI-C" axi_get_temp_static_rw_transaction_write_data_beats_delay = function axi_get_temp_static_rw_transaction_write_data_beats_delay;
    export "DPI-C" axi_set_temp_static_rw_transaction_write_data_beats_delay = function axi_set_temp_static_rw_transaction_write_data_beats_delay;
    export "DPI-C" axi_get_temp_static_rw_transaction_data_valid_delay = function axi_get_temp_static_rw_transaction_data_valid_delay;
    export "DPI-C" axi_set_temp_static_rw_transaction_data_valid_delay = function axi_set_temp_static_rw_transaction_data_valid_delay;
    export "DPI-C" axi_get_temp_static_rw_transaction_data_ready_delay = function axi_get_temp_static_rw_transaction_data_ready_delay;
    export "DPI-C" axi_set_temp_static_rw_transaction_data_ready_delay = function axi_set_temp_static_rw_transaction_data_ready_delay;
    import "DPI-C" context axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog =
    task axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [3:0] burst_length,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] addr_user,
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout axi_rw_e read_or_write,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_valid_delay,
        inout int data_valid_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_response_valid_delay,
        inout int address_ready_delay,
        inout int data_ready_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_response_ready_delay,
        inout bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((4) - 1):0] burst_length,
        inout bit [((8) - 1):0] addr_user,
        inout bit [((8) - 1):0] resp_user,
        inout axi_rw_e read_or_write,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int address_valid_delay,
        inout int write_response_valid_delay,
        inout int address_ready_delay,
        inout int write_response_ready_delay,
        inout bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog =
    task axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_valid_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_ready_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((4) - 1):0] burst_length,
        output bit [((8) - 1):0] addr_user,
        output bit [((8) - 1):0] resp_user,
        output axi_rw_e read_or_write,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        output int address_valid_delay,
        output int write_response_valid_delay,
        output int address_ready_delay,
        output int write_response_ready_delay,
        output bit write_data_with_address,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_AXI_read_addr = function axi_get_temp_static_AXI_read_addr;
    export "DPI-C" axi_set_temp_static_AXI_read_addr = function axi_set_temp_static_AXI_read_addr;
    export "DPI-C" axi_get_temp_static_AXI_read_id = function axi_get_temp_static_AXI_read_id;
    export "DPI-C" axi_set_temp_static_AXI_read_id = function axi_set_temp_static_AXI_read_id;
    export "DPI-C" axi_get_temp_static_AXI_read_data_words = function axi_get_temp_static_AXI_read_data_words;
    export "DPI-C" axi_set_temp_static_AXI_read_data_words = function axi_set_temp_static_AXI_read_data_words;
    export "DPI-C" axi_get_temp_static_AXI_read_resp = function axi_get_temp_static_AXI_read_resp;
    export "DPI-C" axi_set_temp_static_AXI_read_resp = function axi_set_temp_static_AXI_read_resp;
    export "DPI-C" axi_get_temp_static_AXI_read_data_user = function axi_get_temp_static_AXI_read_data_user;
    export "DPI-C" axi_set_temp_static_AXI_read_data_user = function axi_set_temp_static_AXI_read_data_user;
    export "DPI-C" axi_get_temp_static_AXI_read_data_start_time = function axi_get_temp_static_AXI_read_data_start_time;
    export "DPI-C" axi_set_temp_static_AXI_read_data_start_time = function axi_set_temp_static_AXI_read_data_start_time;
    export "DPI-C" axi_get_temp_static_AXI_read_data_end_time = function axi_get_temp_static_AXI_read_data_end_time;
    export "DPI-C" axi_set_temp_static_AXI_read_data_end_time = function axi_set_temp_static_AXI_read_data_end_time;
    import "DPI-C" context axi_AXI_read_ActivatesActivatingActivate_SystemVerilog =
    task axi_AXI_read_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [3:0] burst_length,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] addr_user,
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_to_data_latency,
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((4) - 1):0] burst_length,
        inout bit [((8) - 1):0] addr_user,
        inout int address_to_data_latency,
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_ReceivedReceivingReceive_SystemVerilog =
    task axi_AXI_read_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((4) - 1):0] burst_length,
        output bit [((8) - 1):0] addr_user,
        output int address_to_data_latency,
        output longint addr_start_time,
        output longint addr_end_time,
        output int address_valid_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_AXI_write_addr = function axi_get_temp_static_AXI_write_addr;
    export "DPI-C" axi_set_temp_static_AXI_write_addr = function axi_set_temp_static_AXI_write_addr;
    export "DPI-C" axi_get_temp_static_AXI_write_id = function axi_get_temp_static_AXI_write_id;
    export "DPI-C" axi_set_temp_static_AXI_write_id = function axi_set_temp_static_AXI_write_id;
    export "DPI-C" axi_get_temp_static_AXI_write_data_words = function axi_get_temp_static_AXI_write_data_words;
    export "DPI-C" axi_set_temp_static_AXI_write_data_words = function axi_set_temp_static_AXI_write_data_words;
    export "DPI-C" axi_get_temp_static_AXI_write_write_strobes = function axi_get_temp_static_AXI_write_write_strobes;
    export "DPI-C" axi_set_temp_static_AXI_write_write_strobes = function axi_set_temp_static_AXI_write_write_strobes;
    export "DPI-C" axi_get_temp_static_AXI_write_data_user = function axi_get_temp_static_AXI_write_data_user;
    export "DPI-C" axi_set_temp_static_AXI_write_data_user = function axi_set_temp_static_AXI_write_data_user;
    export "DPI-C" axi_get_temp_static_AXI_write_write_data_beats_delay = function axi_get_temp_static_AXI_write_write_data_beats_delay;
    export "DPI-C" axi_set_temp_static_AXI_write_write_data_beats_delay = function axi_set_temp_static_AXI_write_write_data_beats_delay;
    export "DPI-C" axi_get_temp_static_AXI_write_data_start_time = function axi_get_temp_static_AXI_write_data_start_time;
    export "DPI-C" axi_set_temp_static_AXI_write_data_start_time = function axi_set_temp_static_AXI_write_data_start_time;
    export "DPI-C" axi_get_temp_static_AXI_write_data_end_time = function axi_get_temp_static_AXI_write_data_end_time;
    export "DPI-C" axi_set_temp_static_AXI_write_data_end_time = function axi_set_temp_static_AXI_write_data_end_time;
    import "DPI-C" context axi_AXI_write_ActivatesActivatingActivate_SystemVerilog =
    task axi_AXI_write_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [3:0] burst_length,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout axi_response_e resp,
        inout bit [7:0] addr_user,
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint wr_resp_start_time,
        inout longint wr_resp_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((4) - 1):0] burst_length,
        inout axi_response_e resp,
        inout bit [((8) - 1):0] addr_user,
        inout bit [((8) - 1):0] resp_user,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout longint wr_resp_start_time,
        inout longint wr_resp_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_ReceivedReceivingReceive_SystemVerilog =
    task axi_AXI_write_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((4) - 1):0] burst_length,
        output axi_response_e resp,
        output bit [((8) - 1):0] addr_user,
        output bit [((8) - 1):0] resp_user,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        output longint addr_start_time,
        output longint addr_end_time,
        output longint wr_resp_start_time,
        output longint wr_resp_end_time,
        output int address_valid_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_data_resp_data_words = function axi_get_temp_static_data_resp_data_words;
    export "DPI-C" axi_set_temp_static_data_resp_data_words = function axi_set_temp_static_data_resp_data_words;
    export "DPI-C" axi_get_temp_static_data_resp_write_strobes = function axi_get_temp_static_data_resp_write_strobes;
    export "DPI-C" axi_set_temp_static_data_resp_write_strobes = function axi_set_temp_static_data_resp_write_strobes;
    export "DPI-C" axi_get_temp_static_data_resp_id = function axi_get_temp_static_data_resp_id;
    export "DPI-C" axi_set_temp_static_data_resp_id = function axi_set_temp_static_data_resp_id;
    export "DPI-C" axi_get_temp_static_data_resp_data_user = function axi_get_temp_static_data_resp_data_user;
    export "DPI-C" axi_set_temp_static_data_resp_data_user = function axi_set_temp_static_data_resp_data_user;
    export "DPI-C" axi_get_temp_static_data_resp_write_data_beats_delay = function axi_get_temp_static_data_resp_write_data_beats_delay;
    export "DPI-C" axi_set_temp_static_data_resp_write_data_beats_delay = function axi_set_temp_static_data_resp_write_data_beats_delay;
    export "DPI-C" axi_get_temp_static_data_resp_data_beat_start_time = function axi_get_temp_static_data_resp_data_beat_start_time;
    export "DPI-C" axi_set_temp_static_data_resp_data_beat_start_time = function axi_set_temp_static_data_resp_data_beat_start_time;
    export "DPI-C" axi_get_temp_static_data_resp_data_beat_end_time = function axi_get_temp_static_data_resp_data_beat_end_time;
    export "DPI-C" axi_set_temp_static_data_resp_data_beat_end_time = function axi_set_temp_static_data_resp_data_beat_end_time;
    import "DPI-C" context axi_data_resp_ActivatesActivatingActivate_SystemVerilog =
    task axi_data_resp_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int burst_length,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout axi_response_e resp,
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout longint data_start,
        inout longint data_end,
        inout longint response_start,
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int burst_length,
        inout axi_response_e resp,
        inout bit [((8) - 1):0] resp_user,
        inout longint data_start,
        inout longint data_end,
        inout longint response_start,
        inout longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_ReceivedReceivingReceive_SystemVerilog =
    task axi_data_resp_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output int burst_length,
        output axi_response_e resp,
        output bit [((8) - 1):0] resp_user,
        output longint data_start,
        output longint data_end,
        output longint response_start,
        output longint response_end_time,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_data_burst_data_words = function axi_get_temp_static_read_data_burst_data_words;
    export "DPI-C" axi_set_temp_static_read_data_burst_data_words = function axi_set_temp_static_read_data_burst_data_words;
    export "DPI-C" axi_get_temp_static_read_data_burst_resp = function axi_get_temp_static_read_data_burst_resp;
    export "DPI-C" axi_set_temp_static_read_data_burst_resp = function axi_set_temp_static_read_data_burst_resp;
    export "DPI-C" axi_get_temp_static_read_data_burst_id = function axi_get_temp_static_read_data_burst_id;
    export "DPI-C" axi_set_temp_static_read_data_burst_id = function axi_set_temp_static_read_data_burst_id;
    export "DPI-C" axi_get_temp_static_read_data_burst_data_user = function axi_get_temp_static_read_data_burst_data_user;
    export "DPI-C" axi_set_temp_static_read_data_burst_data_user = function axi_set_temp_static_read_data_burst_data_user;
    export "DPI-C" axi_get_temp_static_read_data_burst_data_start_time = function axi_get_temp_static_read_data_burst_data_start_time;
    export "DPI-C" axi_set_temp_static_read_data_burst_data_start_time = function axi_set_temp_static_read_data_burst_data_start_time;
    export "DPI-C" axi_get_temp_static_read_data_burst_data_end_time = function axi_get_temp_static_read_data_burst_data_end_time;
    export "DPI-C" axi_set_temp_static_read_data_burst_data_end_time = function axi_set_temp_static_read_data_burst_data_end_time;
    import "DPI-C" context axi_read_data_burst_SendSendingSent_SystemVerilog =
    task axi_read_data_burst_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_data_burst_data_words = function axi_get_temp_static_write_data_burst_data_words;
    export "DPI-C" axi_set_temp_static_write_data_burst_data_words = function axi_set_temp_static_write_data_burst_data_words;
    export "DPI-C" axi_get_temp_static_write_data_burst_write_strobes = function axi_get_temp_static_write_data_burst_write_strobes;
    export "DPI-C" axi_set_temp_static_write_data_burst_write_strobes = function axi_set_temp_static_write_data_burst_write_strobes;
    export "DPI-C" axi_get_temp_static_write_data_burst_id = function axi_get_temp_static_write_data_burst_id;
    export "DPI-C" axi_set_temp_static_write_data_burst_id = function axi_set_temp_static_write_data_burst_id;
    export "DPI-C" axi_get_temp_static_write_data_burst_data_user = function axi_get_temp_static_write_data_burst_data_user;
    export "DPI-C" axi_set_temp_static_write_data_burst_data_user = function axi_set_temp_static_write_data_burst_data_user;
    export "DPI-C" axi_get_temp_static_write_data_burst_write_data_beats_delay = function axi_get_temp_static_write_data_burst_write_data_beats_delay;
    export "DPI-C" axi_set_temp_static_write_data_burst_write_data_beats_delay = function axi_set_temp_static_write_data_burst_write_data_beats_delay;
    export "DPI-C" axi_get_temp_static_write_data_burst_data_start_time = function axi_get_temp_static_write_data_burst_data_start_time;
    export "DPI-C" axi_set_temp_static_write_data_burst_data_start_time = function axi_set_temp_static_write_data_burst_data_start_time;
    export "DPI-C" axi_get_temp_static_write_data_burst_data_end_time = function axi_get_temp_static_write_data_burst_data_end_time;
    export "DPI-C" axi_set_temp_static_write_data_burst_data_end_time = function axi_set_temp_static_write_data_burst_data_end_time;
    import "DPI-C" context axi_write_data_burst_SendSendingSent_SystemVerilog =
    task axi_write_data_burst_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int burst_length,
        input int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output int burst_length,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_addr_channel_phase_addr = function axi_get_temp_static_read_addr_channel_phase_addr;
    export "DPI-C" axi_set_temp_static_read_addr_channel_phase_addr = function axi_set_temp_static_read_addr_channel_phase_addr;
    export "DPI-C" axi_get_temp_static_read_addr_channel_phase_id = function axi_get_temp_static_read_addr_channel_phase_id;
    export "DPI-C" axi_set_temp_static_read_addr_channel_phase_id = function axi_set_temp_static_read_addr_channel_phase_id;
    import "DPI-C" context axi_read_addr_channel_phase_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((8) - 1):0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_channel_phase_data = function axi_get_temp_static_read_channel_phase_data;
    export "DPI-C" axi_set_temp_static_read_channel_phase_data = function axi_set_temp_static_read_channel_phase_data;
    export "DPI-C" axi_get_temp_static_read_channel_phase_id = function axi_get_temp_static_read_channel_phase_id;
    export "DPI-C" axi_set_temp_static_read_channel_phase_id = function axi_set_temp_static_read_channel_phase_id;
    import "DPI-C" context axi_read_channel_phase_SendSendingSent_SystemVerilog =
    task axi_read_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input axi_response_e resp,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output axi_response_e resp,
        output bit [((8) - 1):0] data_user,
        output int data_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_addr_channel_phase_addr = function axi_get_temp_static_write_addr_channel_phase_addr;
    export "DPI-C" axi_set_temp_static_write_addr_channel_phase_addr = function axi_set_temp_static_write_addr_channel_phase_addr;
    export "DPI-C" axi_get_temp_static_write_addr_channel_phase_id = function axi_get_temp_static_write_addr_channel_phase_id;
    export "DPI-C" axi_set_temp_static_write_addr_channel_phase_id = function axi_set_temp_static_write_addr_channel_phase_id;
    import "DPI-C" context axi_write_addr_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((8) - 1):0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_channel_phase_data = function axi_get_temp_static_write_channel_phase_data;
    export "DPI-C" axi_set_temp_static_write_channel_phase_data = function axi_set_temp_static_write_channel_phase_data;
    export "DPI-C" axi_get_temp_static_write_channel_phase_write_strobes = function axi_get_temp_static_write_channel_phase_write_strobes;
    export "DPI-C" axi_set_temp_static_write_channel_phase_write_strobes = function axi_set_temp_static_write_channel_phase_write_strobes;
    export "DPI-C" axi_get_temp_static_write_channel_phase_id = function axi_get_temp_static_write_channel_phase_id;
    export "DPI-C" axi_set_temp_static_write_channel_phase_id = function axi_set_temp_static_write_channel_phase_id;
    import "DPI-C" context axi_write_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output bit [((8) - 1):0] data_user,
        output int data_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_resp_channel_phase_id = function axi_get_temp_static_write_resp_channel_phase_id;
    export "DPI-C" axi_set_temp_static_write_resp_channel_phase_id = function axi_set_temp_static_write_resp_channel_phase_id;
    import "DPI-C" context axi_write_resp_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [7:0] resp_user,
        input int write_response_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_resp_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_response_e resp,
        output bit [((8) - 1):0] resp_user,
        output int write_response_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_addr_channel_cycle_addr = function axi_get_temp_static_read_addr_channel_cycle_addr;
    export "DPI-C" axi_set_temp_static_read_addr_channel_cycle_addr = function axi_set_temp_static_read_addr_channel_cycle_addr;
    export "DPI-C" axi_get_temp_static_read_addr_channel_cycle_id = function axi_get_temp_static_read_addr_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_read_addr_channel_cycle_id = function axi_set_temp_static_read_addr_channel_cycle_id;
    import "DPI-C" context axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((8) - 1):0] addr_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_ready_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_channel_cycle_data = function axi_get_temp_static_read_channel_cycle_data;
    export "DPI-C" axi_set_temp_static_read_channel_cycle_data = function axi_set_temp_static_read_channel_cycle_data;
    export "DPI-C" axi_get_temp_static_read_channel_cycle_id = function axi_get_temp_static_read_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_read_channel_cycle_id = function axi_set_temp_static_read_channel_cycle_id;
    import "DPI-C" context axi_read_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_read_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input axi_response_e resp,
        input bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output axi_response_e resp,
        output bit [((8) - 1):0] data_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_ready_SendSendingSent_SystemVerilog =
    task axi_read_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_addr_channel_cycle_addr = function axi_get_temp_static_write_addr_channel_cycle_addr;
    export "DPI-C" axi_set_temp_static_write_addr_channel_cycle_addr = function axi_set_temp_static_write_addr_channel_cycle_addr;
    export "DPI-C" axi_get_temp_static_write_addr_channel_cycle_id = function axi_get_temp_static_write_addr_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_write_addr_channel_cycle_id = function axi_set_temp_static_write_addr_channel_cycle_id;
    import "DPI-C" context axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((8) - 1):0] addr_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_channel_cycle_data = function axi_get_temp_static_write_channel_cycle_data;
    export "DPI-C" axi_set_temp_static_write_channel_cycle_data = function axi_set_temp_static_write_channel_cycle_data;
    export "DPI-C" axi_get_temp_static_write_channel_cycle_strb = function axi_get_temp_static_write_channel_cycle_strb;
    export "DPI-C" axi_set_temp_static_write_channel_cycle_strb = function axi_set_temp_static_write_channel_cycle_strb;
    export "DPI-C" axi_get_temp_static_write_channel_cycle_id = function axi_get_temp_static_write_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_write_channel_cycle_id = function axi_set_temp_static_write_channel_cycle_id;
    import "DPI-C" context axi_write_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output bit [((8) - 1):0] data_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_resp_channel_cycle_id = function axi_get_temp_static_write_resp_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_write_resp_channel_cycle_id = function axi_set_temp_static_write_resp_channel_cycle_id;
    import "DPI-C" context axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [7:0] resp_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_resp_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_response_e resp,
        output bit [((8) - 1):0] resp_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_end_of_timestep_VPI_SystemVerilog =
    task axi_end_of_timestep_VPI_SystemVerilog();
    import "DPI-C" context axi_fn_rd_txn_valid_lanes = function void fn_rd_txn_valid_lanes_C
    (
    );

    import "DPI-C" context axi_fn_get_wdata_phase_info = function void fn_get_wdata_phase_info_C
    (
        input bit wdata_last,
        inout bit waddr_rcvd,
        output bit [3:0] burst_length,
        output int beat_num
    );

    import "DPI-C" context axi_fn_get_wresp_phase_info = function void fn_get_wresp_phase_info_C
    (
    );

    import "DPI-C" context axi_fn_get_rdata_phase_info = function void fn_get_rdata_phase_info_C
    (
        input bit rdata_last,
        output bit [3:0] burst_length,
        output int beat_num
    );

    import "DPI-C" context axi_fn_get_max_os_per_id = function void fn_get_max_os_per_id_C
    (
        output int max_waddr_os,
        output int max_wdata_os
    );

    import "DPI-C" context axi_get_rw_txns_in_prog = function void get_rw_txns_in_prog_C
    (
        output axi_rw_txn_counts_s txn_counts
    );

    import "DPI-C" context axi_fn_add_addr_map_entry = function void fn_add_addr_map_entry_C
    (
        input string region,
        input longint unsigned size
    );

    import "DPI-C" context axi_fn_add_wr_delay = function void fn_add_wr_delay_C
    (
        input string region,
        input bit [17:0] id,
        input int unsigned addr2data,
        input int data2data_DIMS0
    );

    import "DPI-C" context axi_fn_delete_wr_delay = function void fn_delete_wr_delay_C
    (
        input string region,
        input bit [17:0] id
    );

    import "DPI-C" context axi_fn_set_wr_def_delays = function void fn_set_wr_def_delays_C
    (
        input int unsigned min_addr2data,
        input int min_data2data_DIMS0,
        input int unsigned max_addr2data,
        input int max_data2data_DIMS0
    );

    // Waiter task and control
    reg wait_for_control = 0;

    always @(posedge wait_for_control)
    begin
        disable wait_for;
        wait_for_control = 0;
    end

    export "DPI-C" axi_wait_for = task wait_for;

    task wait_for();
        begin
            wait(0 == 1);
        end
    endtask

    // Drive wires (from Cohesive) 
    assign ACLK = internal_ACLK;
    assign ARESETn = internal_ARESETn;
    assign AWVALID = internal_AWVALID;
    assign AWADDR = internal_AWADDR;
    assign AWLEN = internal_AWLEN;
    assign AWSIZE = internal_AWSIZE;
    assign AWBURST = internal_AWBURST;
    assign AWLOCK = internal_AWLOCK;
    assign AWCACHE = internal_AWCACHE;
    assign AWPROT = internal_AWPROT;
    assign AWID = internal_AWID;
    assign AWREADY = internal_AWREADY;
    assign AWUSER = internal_AWUSER;
    assign ARVALID = internal_ARVALID;
    assign ARADDR = internal_ARADDR;
    assign ARLEN = internal_ARLEN;
    assign ARSIZE = internal_ARSIZE;
    assign ARBURST = internal_ARBURST;
    assign ARLOCK = internal_ARLOCK;
    assign ARCACHE = internal_ARCACHE;
    assign ARPROT = internal_ARPROT;
    assign ARID = internal_ARID;
    assign ARREADY = internal_ARREADY;
    assign ARUSER = internal_ARUSER;
    assign RVALID = internal_RVALID;
    assign RLAST = internal_RLAST;
    assign RDATA = internal_RDATA;
    assign RRESP = internal_RRESP;
    assign RID = internal_RID;
    assign RREADY = internal_RREADY;
    assign RUSER = internal_RUSER;
    assign WVALID = internal_WVALID;
    assign WLAST = internal_WLAST;
    assign WDATA = internal_WDATA;
    assign WSTRB = internal_WSTRB;
    assign WID = internal_WID;
    assign WREADY = internal_WREADY;
    assign WUSER = internal_WUSER;
    assign BVALID = internal_BVALID;
    assign BRESP = internal_BRESP;
    assign BID = internal_BID;
    assign BREADY = internal_BREADY;
    assign BUSER = internal_BUSER;
    // Drive wires (from User) 
    assign ACLK = m_ACLK;
    assign ARESETn = m_ARESETn;
    assign AWVALID = m_AWVALID;
    assign AWADDR = m_AWADDR;
    assign AWLEN = m_AWLEN;
    assign AWSIZE = m_AWSIZE;
    assign AWBURST = m_AWBURST;
    assign AWLOCK = m_AWLOCK;
    assign AWCACHE = m_AWCACHE;
    assign AWPROT = m_AWPROT;
    assign AWID = m_AWID;
    assign AWREADY = m_AWREADY;
    assign AWUSER = m_AWUSER;
    assign ARVALID = m_ARVALID;
    assign ARADDR = m_ARADDR;
    assign ARLEN = m_ARLEN;
    assign ARSIZE = m_ARSIZE;
    assign ARBURST = m_ARBURST;
    assign ARLOCK = m_ARLOCK;
    assign ARCACHE = m_ARCACHE;
    assign ARPROT = m_ARPROT;
    assign ARID = m_ARID;
    assign ARREADY = m_ARREADY;
    assign ARUSER = m_ARUSER;
    assign RVALID = m_RVALID;
    assign RLAST = m_RLAST;
    assign RDATA = m_RDATA;
    assign RRESP = m_RRESP;
    assign RID = m_RID;
    assign RREADY = m_RREADY;
    assign RUSER = m_RUSER;
    assign WVALID = m_WVALID;
    assign WLAST = m_WLAST;
    assign WDATA = m_WDATA;
    assign WSTRB = m_WSTRB;
    assign WID = m_WID;
    assign WREADY = m_WREADY;
    assign WUSER = m_WUSER;
    assign BVALID = m_BVALID;
    assign BRESP = m_BRESP;
    assign BID = m_BID;
    assign BREADY = m_BREADY;
    assign BUSER = m_BUSER;

    reg ACLK_changed = 0;
    reg ARESETn_changed = 0;
    reg AWVALID_changed = 0;
    reg AWADDR_changed = 0;
    reg AWLEN_changed = 0;
    reg AWSIZE_changed = 0;
    reg AWBURST_changed = 0;
    reg AWLOCK_changed = 0;
    reg AWCACHE_changed = 0;
    reg AWPROT_changed = 0;
    reg AWID_changed = 0;
    reg AWREADY_changed = 0;
    reg AWUSER_changed = 0;
    reg ARVALID_changed = 0;
    reg ARADDR_changed = 0;
    reg ARLEN_changed = 0;
    reg ARSIZE_changed = 0;
    reg ARBURST_changed = 0;
    reg ARLOCK_changed = 0;
    reg ARCACHE_changed = 0;
    reg ARPROT_changed = 0;
    reg ARID_changed = 0;
    reg ARREADY_changed = 0;
    reg ARUSER_changed = 0;
    reg RVALID_changed = 0;
    reg RLAST_changed = 0;
    reg RDATA_changed = 0;
    reg RRESP_changed = 0;
    reg RID_changed = 0;
    reg RREADY_changed = 0;
    reg RUSER_changed = 0;
    reg WVALID_changed = 0;
    reg WLAST_changed = 0;
    reg WDATA_changed = 0;
    reg WSTRB_changed = 0;
    reg WID_changed = 0;
    reg WREADY_changed = 0;
    reg WUSER_changed = 0;
    reg BVALID_changed = 0;
    reg BRESP_changed = 0;
    reg BID_changed = 0;
    reg BREADY_changed = 0;
    reg BUSER_changed = 0;
    reg config_write_ctrl_to_data_mintime_changed = 0;
    reg config_master_write_delay_changed = 0;
    reg config_enable_all_assertions_changed = 0;
    reg config_enable_assertion_changed = 0;
    reg config_slave_start_addr_changed = 0;
    reg config_slave_end_addr_changed = 0;
    reg config_support_exclusive_access_changed = 0;
    reg config_read_data_reordering_depth_changed = 0;
    reg config_max_transaction_time_factor_changed = 0;
    reg config_timeout_max_data_transfer_changed = 0;
    reg config_burst_timeout_factor_changed = 0;
    reg config_max_latency_AWVALID_assertion_to_AWREADY_changed = 0;
    reg config_max_latency_ARVALID_assertion_to_ARREADY_changed = 0;
    reg config_max_latency_RVALID_assertion_to_RREADY_changed = 0;
    reg config_max_latency_BVALID_assertion_to_BREADY_changed = 0;
    reg config_max_latency_WVALID_assertion_to_WREADY_changed = 0;
    reg config_master_error_position_changed = 0;
    reg config_setup_time_changed = 0;
    reg config_hold_time_changed = 0;
    reg config_max_outstanding_wr_changed = 0;
    reg config_max_outstanding_rd_changed = 0;
    reg config_max_outstanding_rw_changed = 0;
    reg config_is_issuing_changed = 0;

    reg end_of_timestep_control = 0;

    // Start end_of_timestep timer
    initial
    forever
    begin
        wait_end_of_timestep();
    end


    event non_blocking_end_of_timestep_control;

    export "DPI-C" axi_wait_end_of_timestep = task wait_end_of_timestep;

    task wait_end_of_timestep();
        begin
            @(non_blocking_end_of_timestep_control);
            axi_end_of_timestep_VPI_SystemVerilog();
        end
    endtask

    always @( posedge end_of_timestep_control or posedge _check_t0_values )
    begin
        if ( end_of_timestep_control == 1 )
        begin
            ->> non_blocking_end_of_timestep_control;
            end_of_timestep_control = 0;
        end
    end


    // SV wire change monitors

    function automatic void axi_local_set_ACLK_from_SystemVerilog(  );
            axi_set_ACLK_from_SystemVerilog( _interface_ref, ACLK); // DPI call to imported task
        
        axi_propagate_ACLK_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ACLK or posedge _check_t0_values )
    begin
        axi_local_set_ACLK_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARESETn_from_SystemVerilog(  );
            axi_set_ARESETn_from_SystemVerilog( _interface_ref, ARESETn); // DPI call to imported task
        
        axi_propagate_ARESETn_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARESETn or posedge _check_t0_values )
    begin
        axi_local_set_ARESETn_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWVALID_from_SystemVerilog(  );
            axi_set_AWVALID_from_SystemVerilog( _interface_ref, AWVALID); // DPI call to imported task
        
        axi_propagate_AWVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWVALID or posedge _check_t0_values )
    begin
        axi_local_set_AWVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWADDR_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ADDRESS_WIDTH ); _this_dot_1++)
        begin
            axi_set_AWADDR_from_SystemVerilog_index1( _interface_ref, _this_dot_1,AWADDR[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_AWADDR_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWADDR or posedge _check_t0_values )
    begin
        axi_local_set_AWADDR_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWLEN_from_SystemVerilog(  );
            axi_set_AWLEN_from_SystemVerilog( _interface_ref, AWLEN); // DPI call to imported task
        
        axi_propagate_AWLEN_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWLEN or posedge _check_t0_values )
    begin
        axi_local_set_AWLEN_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWSIZE_from_SystemVerilog(  );
            axi_set_AWSIZE_from_SystemVerilog( _interface_ref, AWSIZE); // DPI call to imported task
        
        axi_propagate_AWSIZE_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWSIZE or posedge _check_t0_values )
    begin
        axi_local_set_AWSIZE_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWBURST_from_SystemVerilog(  );
            axi_set_AWBURST_from_SystemVerilog( _interface_ref, AWBURST); // DPI call to imported task
        
        axi_propagate_AWBURST_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWBURST or posedge _check_t0_values )
    begin
        axi_local_set_AWBURST_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWLOCK_from_SystemVerilog(  );
            axi_set_AWLOCK_from_SystemVerilog( _interface_ref, AWLOCK); // DPI call to imported task
        
        axi_propagate_AWLOCK_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWLOCK or posedge _check_t0_values )
    begin
        axi_local_set_AWLOCK_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWCACHE_from_SystemVerilog(  );
            axi_set_AWCACHE_from_SystemVerilog( _interface_ref, AWCACHE); // DPI call to imported task
        
        axi_propagate_AWCACHE_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWCACHE or posedge _check_t0_values )
    begin
        axi_local_set_AWCACHE_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWPROT_from_SystemVerilog(  );
            axi_set_AWPROT_from_SystemVerilog( _interface_ref, AWPROT); // DPI call to imported task
        
        axi_propagate_AWPROT_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWPROT or posedge _check_t0_values )
    begin
        axi_local_set_AWPROT_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_AWID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,AWID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_AWID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWID or posedge _check_t0_values )
    begin
        axi_local_set_AWID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWREADY_from_SystemVerilog(  );
            axi_set_AWREADY_from_SystemVerilog( _interface_ref, AWREADY); // DPI call to imported task
        
        axi_propagate_AWREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWREADY or posedge _check_t0_values )
    begin
        axi_local_set_AWREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWUSER_from_SystemVerilog(  );
            axi_set_AWUSER_from_SystemVerilog( _interface_ref, AWUSER); // DPI call to imported task
        
        axi_propagate_AWUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWUSER or posedge _check_t0_values )
    begin
        axi_local_set_AWUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARVALID_from_SystemVerilog(  );
            axi_set_ARVALID_from_SystemVerilog( _interface_ref, ARVALID); // DPI call to imported task
        
        axi_propagate_ARVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARVALID or posedge _check_t0_values )
    begin
        axi_local_set_ARVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARADDR_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ADDRESS_WIDTH ); _this_dot_1++)
        begin
            axi_set_ARADDR_from_SystemVerilog_index1( _interface_ref, _this_dot_1,ARADDR[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_ARADDR_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARADDR or posedge _check_t0_values )
    begin
        axi_local_set_ARADDR_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARLEN_from_SystemVerilog(  );
            axi_set_ARLEN_from_SystemVerilog( _interface_ref, ARLEN); // DPI call to imported task
        
        axi_propagate_ARLEN_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARLEN or posedge _check_t0_values )
    begin
        axi_local_set_ARLEN_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARSIZE_from_SystemVerilog(  );
            axi_set_ARSIZE_from_SystemVerilog( _interface_ref, ARSIZE); // DPI call to imported task
        
        axi_propagate_ARSIZE_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARSIZE or posedge _check_t0_values )
    begin
        axi_local_set_ARSIZE_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARBURST_from_SystemVerilog(  );
            axi_set_ARBURST_from_SystemVerilog( _interface_ref, ARBURST); // DPI call to imported task
        
        axi_propagate_ARBURST_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARBURST or posedge _check_t0_values )
    begin
        axi_local_set_ARBURST_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARLOCK_from_SystemVerilog(  );
            axi_set_ARLOCK_from_SystemVerilog( _interface_ref, ARLOCK); // DPI call to imported task
        
        axi_propagate_ARLOCK_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARLOCK or posedge _check_t0_values )
    begin
        axi_local_set_ARLOCK_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARCACHE_from_SystemVerilog(  );
            axi_set_ARCACHE_from_SystemVerilog( _interface_ref, ARCACHE); // DPI call to imported task
        
        axi_propagate_ARCACHE_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARCACHE or posedge _check_t0_values )
    begin
        axi_local_set_ARCACHE_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARPROT_from_SystemVerilog(  );
            axi_set_ARPROT_from_SystemVerilog( _interface_ref, ARPROT); // DPI call to imported task
        
        axi_propagate_ARPROT_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARPROT or posedge _check_t0_values )
    begin
        axi_local_set_ARPROT_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_ARID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,ARID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_ARID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARID or posedge _check_t0_values )
    begin
        axi_local_set_ARID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARREADY_from_SystemVerilog(  );
            axi_set_ARREADY_from_SystemVerilog( _interface_ref, ARREADY); // DPI call to imported task
        
        axi_propagate_ARREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARREADY or posedge _check_t0_values )
    begin
        axi_local_set_ARREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARUSER_from_SystemVerilog(  );
            axi_set_ARUSER_from_SystemVerilog( _interface_ref, ARUSER); // DPI call to imported task
        
        axi_propagate_ARUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARUSER or posedge _check_t0_values )
    begin
        axi_local_set_ARUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RVALID_from_SystemVerilog(  );
            axi_set_RVALID_from_SystemVerilog( _interface_ref, RVALID); // DPI call to imported task
        
        axi_propagate_RVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RVALID or posedge _check_t0_values )
    begin
        axi_local_set_RVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RLAST_from_SystemVerilog(  );
            axi_set_RLAST_from_SystemVerilog( _interface_ref, RLAST); // DPI call to imported task
        
        axi_propagate_RLAST_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RLAST or posedge _check_t0_values )
    begin
        axi_local_set_RLAST_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RDATA_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_RDATA_WIDTH ); _this_dot_1++)
        begin
            axi_set_RDATA_from_SystemVerilog_index1( _interface_ref, _this_dot_1,RDATA[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_RDATA_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RDATA or posedge _check_t0_values )
    begin
        axi_local_set_RDATA_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RRESP_from_SystemVerilog(  );
            axi_set_RRESP_from_SystemVerilog( _interface_ref, RRESP); // DPI call to imported task
        
        axi_propagate_RRESP_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RRESP or posedge _check_t0_values )
    begin
        axi_local_set_RRESP_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_RID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,RID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_RID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RID or posedge _check_t0_values )
    begin
        axi_local_set_RID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RREADY_from_SystemVerilog(  );
            axi_set_RREADY_from_SystemVerilog( _interface_ref, RREADY); // DPI call to imported task
        
        axi_propagate_RREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RREADY or posedge _check_t0_values )
    begin
        axi_local_set_RREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RUSER_from_SystemVerilog(  );
            axi_set_RUSER_from_SystemVerilog( _interface_ref, RUSER); // DPI call to imported task
        
        axi_propagate_RUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RUSER or posedge _check_t0_values )
    begin
        axi_local_set_RUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WVALID_from_SystemVerilog(  );
            axi_set_WVALID_from_SystemVerilog( _interface_ref, WVALID); // DPI call to imported task
        
        axi_propagate_WVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WVALID or posedge _check_t0_values )
    begin
        axi_local_set_WVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WLAST_from_SystemVerilog(  );
            axi_set_WLAST_from_SystemVerilog( _interface_ref, WLAST); // DPI call to imported task
        
        axi_propagate_WLAST_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WLAST or posedge _check_t0_values )
    begin
        axi_local_set_WLAST_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WDATA_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_WDATA_WIDTH ); _this_dot_1++)
        begin
            axi_set_WDATA_from_SystemVerilog_index1( _interface_ref, _this_dot_1,WDATA[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_WDATA_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WDATA or posedge _check_t0_values )
    begin
        axi_local_set_WDATA_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WSTRB_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( (AXI_WDATA_WIDTH / 8) ); _this_dot_1++)
        begin
            axi_set_WSTRB_from_SystemVerilog_index1( _interface_ref, _this_dot_1,WSTRB[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_WSTRB_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WSTRB or posedge _check_t0_values )
    begin
        axi_local_set_WSTRB_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_WID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,WID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_WID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WID or posedge _check_t0_values )
    begin
        axi_local_set_WID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WREADY_from_SystemVerilog(  );
            axi_set_WREADY_from_SystemVerilog( _interface_ref, WREADY); // DPI call to imported task
        
        axi_propagate_WREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WREADY or posedge _check_t0_values )
    begin
        axi_local_set_WREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WUSER_from_SystemVerilog(  );
            axi_set_WUSER_from_SystemVerilog( _interface_ref, WUSER); // DPI call to imported task
        
        axi_propagate_WUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WUSER or posedge _check_t0_values )
    begin
        axi_local_set_WUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BVALID_from_SystemVerilog(  );
            axi_set_BVALID_from_SystemVerilog( _interface_ref, BVALID); // DPI call to imported task
        
        axi_propagate_BVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BVALID or posedge _check_t0_values )
    begin
        axi_local_set_BVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BRESP_from_SystemVerilog(  );
            axi_set_BRESP_from_SystemVerilog( _interface_ref, BRESP); // DPI call to imported task
        
        axi_propagate_BRESP_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BRESP or posedge _check_t0_values )
    begin
        axi_local_set_BRESP_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_BID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,BID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_BID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BID or posedge _check_t0_values )
    begin
        axi_local_set_BID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BREADY_from_SystemVerilog(  );
            axi_set_BREADY_from_SystemVerilog( _interface_ref, BREADY); // DPI call to imported task
        
        axi_propagate_BREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BREADY or posedge _check_t0_values )
    begin
        axi_local_set_BREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BUSER_from_SystemVerilog(  );
            axi_set_BUSER_from_SystemVerilog( _interface_ref, BUSER); // DPI call to imported task
        
        axi_propagate_BUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BUSER or posedge _check_t0_values )
    begin
        axi_local_set_BUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end


    // CY wire and variable changed flag monitors

    always @(posedge ACLK_changed or posedge _check_t0_values )
    begin
        while (ACLK_changed == 1'b1)
        begin
            axi_get_ACLK_into_SystemVerilog( _interface_ref, internal_ACLK ); // DPI call to imported task
            ACLK_changed = 1'b0;
            #0  #0 if ( ACLK !== internal_ACLK )
            begin
                axi_local_set_ACLK_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARESETn_changed or posedge _check_t0_values )
    begin
        while (ARESETn_changed == 1'b1)
        begin
            axi_get_ARESETn_into_SystemVerilog( _interface_ref, internal_ARESETn ); // DPI call to imported task
            ARESETn_changed = 1'b0;
            #0  #0 if ( ARESETn !== internal_ARESETn )
            begin
                axi_local_set_ARESETn_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWVALID_changed or posedge _check_t0_values )
    begin
        while (AWVALID_changed == 1'b1)
        begin
            axi_get_AWVALID_into_SystemVerilog( _interface_ref, internal_AWVALID ); // DPI call to imported task
            AWVALID_changed = 1'b0;
            #0  #0 if ( AWVALID !== internal_AWVALID )
            begin
                axi_local_set_AWVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWADDR_changed or posedge _check_t0_values )
    begin
        while (AWADDR_changed == 1'b1)
        begin
            axi_get_AWADDR_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            AWADDR_changed = 1'b0;
            #0  #0 if ( AWADDR !== internal_AWADDR )
            begin
                axi_local_set_AWADDR_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWLEN_changed or posedge _check_t0_values )
    begin
        while (AWLEN_changed == 1'b1)
        begin
            axi_get_AWLEN_into_SystemVerilog( _interface_ref, internal_AWLEN ); // DPI call to imported task
            AWLEN_changed = 1'b0;
            #0  #0 if ( AWLEN !== internal_AWLEN )
            begin
                axi_local_set_AWLEN_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWSIZE_changed or posedge _check_t0_values )
    begin
        while (AWSIZE_changed == 1'b1)
        begin
            axi_get_AWSIZE_into_SystemVerilog( _interface_ref, internal_AWSIZE ); // DPI call to imported task
            AWSIZE_changed = 1'b0;
            #0  #0 if ( AWSIZE !== internal_AWSIZE )
            begin
                axi_local_set_AWSIZE_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWBURST_changed or posedge _check_t0_values )
    begin
        while (AWBURST_changed == 1'b1)
        begin
            axi_get_AWBURST_into_SystemVerilog( _interface_ref, internal_AWBURST ); // DPI call to imported task
            AWBURST_changed = 1'b0;
            #0  #0 if ( AWBURST !== internal_AWBURST )
            begin
                axi_local_set_AWBURST_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWLOCK_changed or posedge _check_t0_values )
    begin
        while (AWLOCK_changed == 1'b1)
        begin
            axi_get_AWLOCK_into_SystemVerilog( _interface_ref, internal_AWLOCK ); // DPI call to imported task
            AWLOCK_changed = 1'b0;
            #0  #0 if ( AWLOCK !== internal_AWLOCK )
            begin
                axi_local_set_AWLOCK_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWCACHE_changed or posedge _check_t0_values )
    begin
        while (AWCACHE_changed == 1'b1)
        begin
            axi_get_AWCACHE_into_SystemVerilog( _interface_ref, internal_AWCACHE ); // DPI call to imported task
            AWCACHE_changed = 1'b0;
            #0  #0 if ( AWCACHE !== internal_AWCACHE )
            begin
                axi_local_set_AWCACHE_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWPROT_changed or posedge _check_t0_values )
    begin
        while (AWPROT_changed == 1'b1)
        begin
            axi_get_AWPROT_into_SystemVerilog( _interface_ref, internal_AWPROT ); // DPI call to imported task
            AWPROT_changed = 1'b0;
            #0  #0 if ( AWPROT !== internal_AWPROT )
            begin
                axi_local_set_AWPROT_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWID_changed or posedge _check_t0_values )
    begin
        while (AWID_changed == 1'b1)
        begin
            axi_get_AWID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            AWID_changed = 1'b0;
            #0  #0 if ( AWID !== internal_AWID )
            begin
                axi_local_set_AWID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWREADY_changed or posedge _check_t0_values )
    begin
        while (AWREADY_changed == 1'b1)
        begin
            axi_get_AWREADY_into_SystemVerilog( _interface_ref, internal_AWREADY ); // DPI call to imported task
            AWREADY_changed = 1'b0;
            #0  #0 if ( AWREADY !== internal_AWREADY )
            begin
                axi_local_set_AWREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWUSER_changed or posedge _check_t0_values )
    begin
        while (AWUSER_changed == 1'b1)
        begin
            axi_get_AWUSER_into_SystemVerilog( _interface_ref, internal_AWUSER ); // DPI call to imported task
            AWUSER_changed = 1'b0;
            #0  #0 if ( AWUSER !== internal_AWUSER )
            begin
                axi_local_set_AWUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARVALID_changed or posedge _check_t0_values )
    begin
        while (ARVALID_changed == 1'b1)
        begin
            axi_get_ARVALID_into_SystemVerilog( _interface_ref, internal_ARVALID ); // DPI call to imported task
            ARVALID_changed = 1'b0;
            #0  #0 if ( ARVALID !== internal_ARVALID )
            begin
                axi_local_set_ARVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARADDR_changed or posedge _check_t0_values )
    begin
        while (ARADDR_changed == 1'b1)
        begin
            axi_get_ARADDR_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            ARADDR_changed = 1'b0;
            #0  #0 if ( ARADDR !== internal_ARADDR )
            begin
                axi_local_set_ARADDR_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARLEN_changed or posedge _check_t0_values )
    begin
        while (ARLEN_changed == 1'b1)
        begin
            axi_get_ARLEN_into_SystemVerilog( _interface_ref, internal_ARLEN ); // DPI call to imported task
            ARLEN_changed = 1'b0;
            #0  #0 if ( ARLEN !== internal_ARLEN )
            begin
                axi_local_set_ARLEN_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARSIZE_changed or posedge _check_t0_values )
    begin
        while (ARSIZE_changed == 1'b1)
        begin
            axi_get_ARSIZE_into_SystemVerilog( _interface_ref, internal_ARSIZE ); // DPI call to imported task
            ARSIZE_changed = 1'b0;
            #0  #0 if ( ARSIZE !== internal_ARSIZE )
            begin
                axi_local_set_ARSIZE_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARBURST_changed or posedge _check_t0_values )
    begin
        while (ARBURST_changed == 1'b1)
        begin
            axi_get_ARBURST_into_SystemVerilog( _interface_ref, internal_ARBURST ); // DPI call to imported task
            ARBURST_changed = 1'b0;
            #0  #0 if ( ARBURST !== internal_ARBURST )
            begin
                axi_local_set_ARBURST_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARLOCK_changed or posedge _check_t0_values )
    begin
        while (ARLOCK_changed == 1'b1)
        begin
            axi_get_ARLOCK_into_SystemVerilog( _interface_ref, internal_ARLOCK ); // DPI call to imported task
            ARLOCK_changed = 1'b0;
            #0  #0 if ( ARLOCK !== internal_ARLOCK )
            begin
                axi_local_set_ARLOCK_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARCACHE_changed or posedge _check_t0_values )
    begin
        while (ARCACHE_changed == 1'b1)
        begin
            axi_get_ARCACHE_into_SystemVerilog( _interface_ref, internal_ARCACHE ); // DPI call to imported task
            ARCACHE_changed = 1'b0;
            #0  #0 if ( ARCACHE !== internal_ARCACHE )
            begin
                axi_local_set_ARCACHE_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARPROT_changed or posedge _check_t0_values )
    begin
        while (ARPROT_changed == 1'b1)
        begin
            axi_get_ARPROT_into_SystemVerilog( _interface_ref, internal_ARPROT ); // DPI call to imported task
            ARPROT_changed = 1'b0;
            #0  #0 if ( ARPROT !== internal_ARPROT )
            begin
                axi_local_set_ARPROT_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARID_changed or posedge _check_t0_values )
    begin
        while (ARID_changed == 1'b1)
        begin
            axi_get_ARID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            ARID_changed = 1'b0;
            #0  #0 if ( ARID !== internal_ARID )
            begin
                axi_local_set_ARID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARREADY_changed or posedge _check_t0_values )
    begin
        while (ARREADY_changed == 1'b1)
        begin
            axi_get_ARREADY_into_SystemVerilog( _interface_ref, internal_ARREADY ); // DPI call to imported task
            ARREADY_changed = 1'b0;
            #0  #0 if ( ARREADY !== internal_ARREADY )
            begin
                axi_local_set_ARREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARUSER_changed or posedge _check_t0_values )
    begin
        while (ARUSER_changed == 1'b1)
        begin
            axi_get_ARUSER_into_SystemVerilog( _interface_ref, internal_ARUSER ); // DPI call to imported task
            ARUSER_changed = 1'b0;
            #0  #0 if ( ARUSER !== internal_ARUSER )
            begin
                axi_local_set_ARUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RVALID_changed or posedge _check_t0_values )
    begin
        while (RVALID_changed == 1'b1)
        begin
            axi_get_RVALID_into_SystemVerilog( _interface_ref, internal_RVALID ); // DPI call to imported task
            RVALID_changed = 1'b0;
            #0  #0 if ( RVALID !== internal_RVALID )
            begin
                axi_local_set_RVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RLAST_changed or posedge _check_t0_values )
    begin
        while (RLAST_changed == 1'b1)
        begin
            axi_get_RLAST_into_SystemVerilog( _interface_ref, internal_RLAST ); // DPI call to imported task
            RLAST_changed = 1'b0;
            #0  #0 if ( RLAST !== internal_RLAST )
            begin
                axi_local_set_RLAST_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RDATA_changed or posedge _check_t0_values )
    begin
        while (RDATA_changed == 1'b1)
        begin
            axi_get_RDATA_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            RDATA_changed = 1'b0;
            #0  #0 if ( RDATA !== internal_RDATA )
            begin
                axi_local_set_RDATA_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RRESP_changed or posedge _check_t0_values )
    begin
        while (RRESP_changed == 1'b1)
        begin
            axi_get_RRESP_into_SystemVerilog( _interface_ref, internal_RRESP ); // DPI call to imported task
            RRESP_changed = 1'b0;
            #0  #0 if ( RRESP !== internal_RRESP )
            begin
                axi_local_set_RRESP_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RID_changed or posedge _check_t0_values )
    begin
        while (RID_changed == 1'b1)
        begin
            axi_get_RID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            RID_changed = 1'b0;
            #0  #0 if ( RID !== internal_RID )
            begin
                axi_local_set_RID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RREADY_changed or posedge _check_t0_values )
    begin
        while (RREADY_changed == 1'b1)
        begin
            axi_get_RREADY_into_SystemVerilog( _interface_ref, internal_RREADY ); // DPI call to imported task
            RREADY_changed = 1'b0;
            #0  #0 if ( RREADY !== internal_RREADY )
            begin
                axi_local_set_RREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RUSER_changed or posedge _check_t0_values )
    begin
        while (RUSER_changed == 1'b1)
        begin
            axi_get_RUSER_into_SystemVerilog( _interface_ref, internal_RUSER ); // DPI call to imported task
            RUSER_changed = 1'b0;
            #0  #0 if ( RUSER !== internal_RUSER )
            begin
                axi_local_set_RUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WVALID_changed or posedge _check_t0_values )
    begin
        while (WVALID_changed == 1'b1)
        begin
            axi_get_WVALID_into_SystemVerilog( _interface_ref, internal_WVALID ); // DPI call to imported task
            WVALID_changed = 1'b0;
            #0  #0 if ( WVALID !== internal_WVALID )
            begin
                axi_local_set_WVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WLAST_changed or posedge _check_t0_values )
    begin
        while (WLAST_changed == 1'b1)
        begin
            axi_get_WLAST_into_SystemVerilog( _interface_ref, internal_WLAST ); // DPI call to imported task
            WLAST_changed = 1'b0;
            #0  #0 if ( WLAST !== internal_WLAST )
            begin
                axi_local_set_WLAST_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WDATA_changed or posedge _check_t0_values )
    begin
        while (WDATA_changed == 1'b1)
        begin
            axi_get_WDATA_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            WDATA_changed = 1'b0;
            #0  #0 if ( WDATA !== internal_WDATA )
            begin
                axi_local_set_WDATA_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WSTRB_changed or posedge _check_t0_values )
    begin
        while (WSTRB_changed == 1'b1)
        begin
            axi_get_WSTRB_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            WSTRB_changed = 1'b0;
            #0  #0 if ( WSTRB !== internal_WSTRB )
            begin
                axi_local_set_WSTRB_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WID_changed or posedge _check_t0_values )
    begin
        while (WID_changed == 1'b1)
        begin
            axi_get_WID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            WID_changed = 1'b0;
            #0  #0 if ( WID !== internal_WID )
            begin
                axi_local_set_WID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WREADY_changed or posedge _check_t0_values )
    begin
        while (WREADY_changed == 1'b1)
        begin
            axi_get_WREADY_into_SystemVerilog( _interface_ref, internal_WREADY ); // DPI call to imported task
            WREADY_changed = 1'b0;
            #0  #0 if ( WREADY !== internal_WREADY )
            begin
                axi_local_set_WREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WUSER_changed or posedge _check_t0_values )
    begin
        while (WUSER_changed == 1'b1)
        begin
            axi_get_WUSER_into_SystemVerilog( _interface_ref, internal_WUSER ); // DPI call to imported task
            WUSER_changed = 1'b0;
            #0  #0 if ( WUSER !== internal_WUSER )
            begin
                axi_local_set_WUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BVALID_changed or posedge _check_t0_values )
    begin
        while (BVALID_changed == 1'b1)
        begin
            axi_get_BVALID_into_SystemVerilog( _interface_ref, internal_BVALID ); // DPI call to imported task
            BVALID_changed = 1'b0;
            #0  #0 if ( BVALID !== internal_BVALID )
            begin
                axi_local_set_BVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BRESP_changed or posedge _check_t0_values )
    begin
        while (BRESP_changed == 1'b1)
        begin
            axi_get_BRESP_into_SystemVerilog( _interface_ref, internal_BRESP ); // DPI call to imported task
            BRESP_changed = 1'b0;
            #0  #0 if ( BRESP !== internal_BRESP )
            begin
                axi_local_set_BRESP_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BID_changed or posedge _check_t0_values )
    begin
        while (BID_changed == 1'b1)
        begin
            axi_get_BID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            BID_changed = 1'b0;
            #0  #0 if ( BID !== internal_BID )
            begin
                axi_local_set_BID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BREADY_changed or posedge _check_t0_values )
    begin
        while (BREADY_changed == 1'b1)
        begin
            axi_get_BREADY_into_SystemVerilog( _interface_ref, internal_BREADY ); // DPI call to imported task
            BREADY_changed = 1'b0;
            #0  #0 if ( BREADY !== internal_BREADY )
            begin
                axi_local_set_BREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BUSER_changed or posedge _check_t0_values )
    begin
        while (BUSER_changed == 1'b1)
        begin
            axi_get_BUSER_into_SystemVerilog( _interface_ref, internal_BUSER ); // DPI call to imported task
            BUSER_changed = 1'b0;
            #0  #0 if ( BUSER !== internal_BUSER )
            begin
                axi_local_set_BUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge config_write_ctrl_to_data_mintime_changed or posedge _check_t0_values )
    begin
        if (config_write_ctrl_to_data_mintime_changed == 1'b1)
        begin
            axi_get_config_write_ctrl_to_data_mintime_into_SystemVerilog( _interface_ref, config_write_ctrl_to_data_mintime ); // DPI call to imported task
            config_write_ctrl_to_data_mintime_changed = 1'b0;
        end
    end

    always @(posedge config_master_write_delay_changed or posedge _check_t0_values )
    begin
        if (config_master_write_delay_changed == 1'b1)
        begin
            axi_get_config_master_write_delay_into_SystemVerilog( _interface_ref, config_master_write_delay ); // DPI call to imported task
            config_master_write_delay_changed = 1'b0;
        end
    end

    always @(posedge config_enable_all_assertions_changed or posedge _check_t0_values )
    begin
        if (config_enable_all_assertions_changed == 1'b1)
        begin
            axi_get_config_enable_all_assertions_into_SystemVerilog( _interface_ref, config_enable_all_assertions ); // DPI call to imported task
            config_enable_all_assertions_changed = 1'b0;
        end
    end

    always @(posedge config_enable_assertion_changed or posedge _check_t0_values )
    begin
        if (config_enable_assertion_changed == 1'b1)
        begin
            axi_get_config_enable_assertion_into_SystemVerilog( _interface_ref, config_enable_assertion ); // DPI call to imported task
            config_enable_assertion_changed = 1'b0;
        end
    end

    always @(posedge config_slave_start_addr_changed or posedge _check_t0_values )
    begin
        if (config_slave_start_addr_changed == 1'b1)
        begin
            axi_get_config_slave_start_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            config_slave_start_addr_changed = 1'b0;
        end
    end

    always @(posedge config_slave_end_addr_changed or posedge _check_t0_values )
    begin
        if (config_slave_end_addr_changed == 1'b1)
        begin
            axi_get_config_slave_end_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            config_slave_end_addr_changed = 1'b0;
        end
    end

    always @(posedge config_support_exclusive_access_changed or posedge _check_t0_values )
    begin
        if (config_support_exclusive_access_changed == 1'b1)
        begin
            axi_get_config_support_exclusive_access_into_SystemVerilog( _interface_ref, config_support_exclusive_access ); // DPI call to imported task
            config_support_exclusive_access_changed = 1'b0;
        end
    end

    always @(posedge config_read_data_reordering_depth_changed or posedge _check_t0_values )
    begin
        if (config_read_data_reordering_depth_changed == 1'b1)
        begin
            axi_get_config_read_data_reordering_depth_into_SystemVerilog( _interface_ref, config_read_data_reordering_depth ); // DPI call to imported task
            config_read_data_reordering_depth_changed = 1'b0;
        end
    end

    always @(posedge config_max_transaction_time_factor_changed or posedge _check_t0_values )
    begin
        if (config_max_transaction_time_factor_changed == 1'b1)
        begin
            axi_get_config_max_transaction_time_factor_into_SystemVerilog( _interface_ref, config_max_transaction_time_factor ); // DPI call to imported task
            config_max_transaction_time_factor_changed = 1'b0;
        end
    end

    always @(posedge config_timeout_max_data_transfer_changed or posedge _check_t0_values )
    begin
        if (config_timeout_max_data_transfer_changed == 1'b1)
        begin
            axi_get_config_timeout_max_data_transfer_into_SystemVerilog( _interface_ref, config_timeout_max_data_transfer ); // DPI call to imported task
            config_timeout_max_data_transfer_changed = 1'b0;
        end
    end

    always @(posedge config_burst_timeout_factor_changed or posedge _check_t0_values )
    begin
        if (config_burst_timeout_factor_changed == 1'b1)
        begin
            axi_get_config_burst_timeout_factor_into_SystemVerilog( _interface_ref, config_burst_timeout_factor ); // DPI call to imported task
            config_burst_timeout_factor_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_AWVALID_assertion_to_AWREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_AWVALID_assertion_to_AWREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_AWVALID_assertion_to_AWREADY_into_SystemVerilog( _interface_ref, config_max_latency_AWVALID_assertion_to_AWREADY ); // DPI call to imported task
            config_max_latency_AWVALID_assertion_to_AWREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_ARVALID_assertion_to_ARREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_ARVALID_assertion_to_ARREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_ARVALID_assertion_to_ARREADY_into_SystemVerilog( _interface_ref, config_max_latency_ARVALID_assertion_to_ARREADY ); // DPI call to imported task
            config_max_latency_ARVALID_assertion_to_ARREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_RVALID_assertion_to_RREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_RVALID_assertion_to_RREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_RVALID_assertion_to_RREADY_into_SystemVerilog( _interface_ref, config_max_latency_RVALID_assertion_to_RREADY ); // DPI call to imported task
            config_max_latency_RVALID_assertion_to_RREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_BVALID_assertion_to_BREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_BVALID_assertion_to_BREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_BVALID_assertion_to_BREADY_into_SystemVerilog( _interface_ref, config_max_latency_BVALID_assertion_to_BREADY ); // DPI call to imported task
            config_max_latency_BVALID_assertion_to_BREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_WVALID_assertion_to_WREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_WVALID_assertion_to_WREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_WVALID_assertion_to_WREADY_into_SystemVerilog( _interface_ref, config_max_latency_WVALID_assertion_to_WREADY ); // DPI call to imported task
            config_max_latency_WVALID_assertion_to_WREADY_changed = 1'b0;
        end
    end

    always @(posedge config_master_error_position_changed or posedge _check_t0_values )
    begin
        if (config_master_error_position_changed == 1'b1)
        begin
            axi_get_config_master_error_position_into_SystemVerilog( _interface_ref, config_master_error_position ); // DPI call to imported task
            config_master_error_position_changed = 1'b0;
        end
    end

    always @(posedge config_setup_time_changed or posedge _check_t0_values )
    begin
        if (config_setup_time_changed == 1'b1)
        begin
            axi_get_config_setup_time_into_SystemVerilog( _interface_ref, config_setup_time ); // DPI call to imported task
            config_setup_time_changed = 1'b0;
        end
    end

    always @(posedge config_hold_time_changed or posedge _check_t0_values )
    begin
        if (config_hold_time_changed == 1'b1)
        begin
            axi_get_config_hold_time_into_SystemVerilog( _interface_ref, config_hold_time ); // DPI call to imported task
            config_hold_time_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_wr_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_wr_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_wr_into_SystemVerilog( _interface_ref, config_max_outstanding_wr ); // DPI call to imported task
            config_max_outstanding_wr_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_rd_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_rd_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_rd_into_SystemVerilog( _interface_ref, config_max_outstanding_rd ); // DPI call to imported task
            config_max_outstanding_rd_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_rw_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_rw_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_rw_into_SystemVerilog( _interface_ref, config_max_outstanding_rw ); // DPI call to imported task
            config_max_outstanding_rw_changed = 1'b0;
        end
    end

    always @(posedge config_is_issuing_changed or posedge _check_t0_values )
    begin
        if (config_is_issuing_changed == 1'b1)
        begin
            axi_get_config_is_issuing_into_SystemVerilog( _interface_ref, config_is_issuing ); // DPI call to imported task
            config_is_issuing_changed = 1'b0;
        end
    end


    //--------------------------------------------------------------------------------
    // Task which blocks and outputs an error if the interface has not initialized properly
    //--------------------------------------------------------------------------------

    task _initialized();
        if (_interface_ref == 0)
        begin
            $display("Error: %m - Questa Verification IP failed to initialise. Please check questa_mvc.log for details");
            wait(_interface_ref!=0);
        end
    endtask

endinterface

`endif // INCA
`ifdef VCS
// *****************************************************************************
//
// Copyright 2007-2016 Mentor Graphics Corporation
// All Rights Reserved.
//
// THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE PROPERTY OF
// MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS.
//
// *****************************************************************************
// SystemVerilog           Version: 20160107
// *****************************************************************************

import QUESTA_MVC::questa_mvc_reporter;
import QUESTA_MVC::questa_mvc_item_comms_semantic;
import QUESTA_MVC::questa_mvc_edge;
import QUESTA_MVC::QUESTA_MVC_POSEDGE;
import QUESTA_MVC::QUESTA_MVC_NEGEDGE;
import QUESTA_MVC::QUESTA_MVC_ANYEDGE;
import QUESTA_MVC::QUESTA_MVC_0_TO_1_EDGE;
import QUESTA_MVC::QUESTA_MVC_1_TO_0_EDGE;


(* cy_so="libaxi_IN_SystemVerilog_MTI_full" *)
(* on_lib_load="axi_IN_SystemVerilog_load" *)

interface mgc_common_axi #(int AXI_ADDRESS_WIDTH = 64, int AXI_RDATA_WIDTH = 1024, int AXI_WDATA_WIDTH = 1024, int AXI_ID_WIDTH = 18)
    (input wire iACLK, input wire iARESETn);

    //-------------------------------------------------------------------------
    //
    // Group: AXI Signals
    //
    //-------------------------------------------------------------------------



    //-------------------------------------------------------------------------
    // Private wires
    //-------------------------------------------------------------------------
    wire ACLK;
    wire ARESETn;
    wire AWVALID;
    wire [((AXI_ADDRESS_WIDTH) - 1):0]  AWADDR;
    wire [3:0] AWLEN;
    wire [2:0] AWSIZE;
    wire [1:0] AWBURST;
    wire [1:0] AWLOCK;
    wire [3:0] AWCACHE;
    wire [2:0] AWPROT;
    wire [((AXI_ID_WIDTH) - 1):0]  AWID;
    wire AWREADY;
    wire [7:0] AWUSER;
    wire ARVALID;
    wire [((AXI_ADDRESS_WIDTH) - 1):0]  ARADDR;
    wire [3:0] ARLEN;
    wire [2:0] ARSIZE;
    wire [1:0] ARBURST;
    wire [1:0] ARLOCK;
    wire [3:0] ARCACHE;
    wire [2:0] ARPROT;
    wire [((AXI_ID_WIDTH) - 1):0]  ARID;
    wire ARREADY;
    wire [7:0] ARUSER;
    wire RVALID;
    wire RLAST;
    wire [((AXI_RDATA_WIDTH) - 1):0]  RDATA;
    wire [1:0] RRESP;
    wire [((AXI_ID_WIDTH) - 1):0]  RID;
    wire RREADY;
    wire [7:0] RUSER;
    wire WVALID;
    wire WLAST;
    wire [((AXI_WDATA_WIDTH) - 1):0]  WDATA;
    wire [(((AXI_WDATA_WIDTH / 8)) - 1):0]  WSTRB;
    wire [((AXI_ID_WIDTH) - 1):0]  WID;
    wire WREADY;
    wire [7:0] WUSER;
    wire BVALID;
    wire [1:0] BRESP;
    wire [((AXI_ID_WIDTH) - 1):0]  BID;
    wire BREADY;
    wire [7:0] BUSER;



    // Propagate global signals onto interface wires
    assign ACLK = iACLK;
    assign ARESETn = iARESETn;

    // Variable: config_write_ctrl_to_data_mintime
    //
    // 
    // Sets the delay from start of address phase to start of data phase in a write 
    // transaction (in terms of ACLK).
    // 
    // Default: 1 
    // 
    // This configuration variable has been deprecated and is maintained 
    // for backward compatibility. However, you can use ~write_address_to_data_delay~ 
    // configuration variable to control the delay between a write address phase 
    // and a write data phase.
    // 
    //
    int unsigned config_write_ctrl_to_data_mintime;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Enables
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_enable_all_assertions
    //
    // 
    // Enables all protocol assertions. 
    // 
    // Default: 1
    // 
    //
    // mentor configurator specification name "Enable all protocol assertions"
    bit config_enable_all_assertions;

    // Variable: config_enable_assertion
    //
    // 
    // Enables individual protocol assertion.
    // This variable controls whether specific assertion within QVIP (of type <axi_assertion_e>) is enabled or disabled.
    // Individual assertion can be disabled as follows:-
    // //-----------------------------------------------------------------------
    // // < BFM interface>.set_config_enable_assertion_index1(<name of assertion>,1'b0);
    // //-----------------------------------------------------------------------
    // 
    // For example, the assertion AXI_READ_DATA_UNKN is disabled as follows:
    // <bfm>.set_config_enable_assertion_index1(AXI_READ_DATA_UNKN, 1'b0); 
    // 
    // Here bfm is the AXI interface instance name for which the assertion to be disabled. 
    // 
    // Default: All assertions are enabled
    //   
    // 
    //
    // mentor configurator specification name "Enable individual protocol assertion"
    bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Slave behavior control
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_support_exclusive_access
    //
    // 
    // Enables exclusive transactions support for slave.
    // If disabled, every exclusive read/write returns an OKAY response,
    // and exclusive write updates memory. 
    // 
    // Default: 1  
    // 
    //
    // mentor configurator specification name "Enable exclusive transaction support"
    bit config_support_exclusive_access;

    // Variable: config_read_data_reordering_depth
    //
    // 
    // Sets the maximum number of different read transaction addresses for which read 
    // data(response) can be sent in any order from slave. 
    // 
    // Default: 2 ** AXI_ID_WIDTH
    // 
    //
    // mentor configurator specification name "Read data reordering depth"
    int unsigned config_read_data_reordering_depth;

    // 
    // //-----------------------------------------------------------------------------
    // Group: Timeout control
    // //-----------------------------------------------------------------------------
    // 


    // Variable: config_max_transaction_time_factor
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) for any complete read or write transaction, which
    // includes time period for all individual phases of transaction. 
    // 
    // Default: 100000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout for complete read/write transaction"
    int unsigned config_max_transaction_time_factor;

    // Variable: config_timeout_max_data_transfer
    //
    //  
    // Sets maximum number of write data beats in a write data burst. 
    // 
    // Default: 1024  
    // 
    //
    // mentor configurator specification name "Maximum number of data beats in a write data burst"
    int config_timeout_max_data_transfer;

    // Variable: config_burst_timeout_factor
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) between individual phases of a transaction. 
    // 
    // Default: 10000 clock cycles 
    // 
    //
    // mentor configurator specification name "Burst timeout between individual phases of a transaction"
    int unsigned config_burst_timeout_factor;

    // Variable: config_max_latency_AWVALID_assertion_to_AWREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of AWVALID to assertion of AWREADY.
    // An error message AXI_AWREADY_NOT_ASSERTED_AFTER_AWVALID is generated if AWREADY is not asserted
    // after assertion of AWVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from AWVALID to AWREADY assertion"
    int unsigned config_max_latency_AWVALID_assertion_to_AWREADY;

    // Variable: config_max_latency_ARVALID_assertion_to_ARREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of ARVALID to assertion of ARREADY.
    // An error message AXI_ARREADY_NOT_ASSERTED_AFTER_ARVALID is generated if ARREADY is not asserted
    // after assertion of ARVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from ARVALID to ARREADY assertion"
    int unsigned config_max_latency_ARVALID_assertion_to_ARREADY;

    // Variable: config_max_latency_RVALID_assertion_to_RREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of RVALID to assertion of RREADY.
    // An error message AXI_RREADY_NOT_ASSERTED_AFTER_RVALID is generated if RREADY is not asserted
    // after assertion of RVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from RVALID to RREADY assertion"
    int unsigned config_max_latency_RVALID_assertion_to_RREADY;

    // Variable: config_max_latency_BVALID_assertion_to_BREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of BVALID to assertion of BREADY.
    // An error message AXI_BREADY_NOT_ASSERTED_AFTER_BVALID is generated if BREADY is not asserted
    // after assertion of BVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from BVALID to BREADY assertion"
    int unsigned config_max_latency_BVALID_assertion_to_BREADY;

    // Variable: config_max_latency_WVALID_assertion_to_WREADY
    //
    //  
    // Sets maximum timeout period (in terms of ACLK) from assertion of WVALID to assertion of WREADY.
    // An error message AXI_WREADY_NOT_ASSERTED_AFTER_WVALID is generated if WREADY is not asserted
    // after assertion of WVALID within this period. 
    // 
    // Default: 10000 clock cycles
    // 
    //
    // mentor configurator specification name "Timeout from WVALID to WREADY assertion"
    int unsigned config_max_latency_WVALID_assertion_to_WREADY;

    // Variable: config_setup_time
    //
    // 
    // Sets number of simulation time units from the setup time to the active 
    // clock edge of ACLK. The setup time will always be less than the time period
    // of the clock. 
    // 
    // Default: 0
    // 
    //
    // Note - This configuration variable is used in an expression involving time precision.
    //        To ensure its value is correct, use questa_mvc_sv_convert_to_precision API of QUESTA_MVC package.
    //
    int config_setup_time;

    // Variable: config_hold_time
    //
    // 
    // Sets number of simulation time units from the hold time to the active 
    // clock edge of ACLK. 
    // 
    // Default: 0
    // 
    //
    // Note - This configuration variable is used in an expression involving time precision.
    //        To ensure its value is correct, use questa_mvc_sv_convert_to_precision API of QUESTA_MVC package.
    //
    int config_hold_time;

    // Variable: config_max_outstanding_wr
    //
    // Configures maximum possible outstanding Write transactions
    //
    int config_max_outstanding_wr;

    // Variable: config_max_outstanding_rd
    //
    // Configures maximum possible outstanding Read transactions
    //
    int config_max_outstanding_rd;

    // Variable: config_max_outstanding_rw
    //
    // Configures maximum possible outstanding Combined (Read and Write) transactions
    //
    int config_max_outstanding_rw;

    // Variable: config_is_issuing
    //
    // Enables Master component to use "config_max_outstanding_wr/config_max_outstanding_rd/config_max_outstanding_rw" variables for transaction issuing capability when set to true
    //
    bit config_is_issuing;


    //-------------------------------------------------------------------------
    // Deprecated variables - writing to these variables will cause a warning to be issued.
    //-------------------------------------------------------------------------
    bit config_master_write_delay;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr;
    axi_error_e config_master_error_position;
    //------------------------------------------------------------------------------
    // Group:- Interface ends
    //------------------------------------------------------------------------------
    //
    longint axi_master_end;


    // Function:- get_axi_master_end
    //
    // Returns a handle to the <master> end of this instance of the <axi> interface.

    function longint get_axi_master_end();
        return axi_master_end;
    endfunction

    longint axi_slave_end;


    // Function:- get_axi_slave_end
    //
    // Returns a handle to the <slave> end of this instance of the <axi> interface.

    function longint get_axi_slave_end();
        return axi_slave_end;
    endfunction

    longint axi_clock_source_end;


    // Function:- get_axi_clock_source_end
    //
    // Returns a handle to the <clock_source> end of this instance of the <axi> interface.

    function longint get_axi_clock_source_end();
        return axi_clock_source_end;
    endfunction

    longint axi_reset_source_end;


    // Function:- get_axi_reset_source_end
    //
    // Returns a handle to the <reset_source> end of this instance of the <axi> interface.

    function longint get_axi_reset_source_end();
        return axi_reset_source_end;
    endfunction

    longint axi__monitor_end;


    // Function:- get_axi__monitor_end
    //
    // Returns a handle to the <_monitor> end of this instance of the <axi> interface.

    function longint get_axi__monitor_end();
        return axi__monitor_end;
    endfunction


    // Group:- Abstraction Levels
    // 
    // These functions are used set or get the abstraction levels of an interface end.
    // See <Abstraction Levels of Interface Ends> for more details on the meaning of
    // TLM or WLM connected and the valid combinations.


    //-------------------------------------------------------------------------
    // Function:- axi_set_master_abstraction_level
    //
    //     Function to set whether the <master> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_master_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_master_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_master_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <master> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_master_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_master_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_slave_abstraction_level
    //
    //     Function to set whether the <slave> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_slave_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_slave_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_slave_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <slave> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_slave_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_slave_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_clock_source_abstraction_level
    //
    //     Function to set whether the <clock_source> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_clock_source_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_clock_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_clock_source_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <clock_source> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_clock_source_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_clock_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_set_reset_source_abstraction_level
    //
    //     Function to set whether the <reset_source> end of the interface is WLM
    //     or TLM connected. See <Abstraction Levels of Interface Ends> for a
    //     description of abstraction levels, how they affect the behaviour of the
    //     QVIP, and guidelines for setting them.
    //
    // Arguments:
    //    wire_level - Set to 1 to be WLM connected.
    //    TLM_level -  Set to 1 to be TLM connected.
    //
    function void axi_set_reset_source_abstraction_level
    (
        input bit          wire_level,
        input bit          TLM_level
    );
        axi_set_reset_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- axi_get_reset_source_abstraction_level
    //
    //     Function to return the Abstraction level setting for the <reset_source> end.
    //     See <Abstraction Levels of Interface Ends> for a description of abstraction
    //     levels and how they affect the behaviour of the Questa Verification IP.
    //
    // Arguments:
    //
    //    wire_level - Value = 1 if this end is WLM connected.
    //    TLM_level -  Value = 1 if this end is TLM connected.
    //------------------------------------------------------------------------------
    function void axi_get_reset_source_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
        axi_get_reset_source_end_abstraction_level( wire_level, TLM_level );
    endfunction

    import "DPI-C" context function longint axi_initialise_SystemVerilog
    (
        int    usage_code,
        string iface_version,
        output longint master_end,
        output longint slave_end,
        output longint clock_source_end,
        output longint reset_source_end,
        output longint _monitor_end,
        input int AXI_ADDRESS_WIDTH,
        input int AXI_RDATA_WIDTH,
        input int AXI_WDATA_WIDTH,
        input int AXI_ID_WIDTH
    );

    `ifndef MVC_axi_VERSION
    `define MVC_axi_VERSION ""
    `endif
    // Handle to the linkage
    (* elab_init *) longint _interface_ref =
                                axi_initialise_SystemVerilog
                                (
                                    18102076,
                                    `MVC_axi_VERSION,
                                    axi_master_end,
                                    axi_slave_end,
                                    axi_clock_source_end,
                                    axi_reset_source_end,
                                    axi__monitor_end,
                                    AXI_ADDRESS_WIDTH,
                                    AXI_RDATA_WIDTH,
                                    AXI_WDATA_WIDTH,
                                    AXI_ID_WIDTH
                                ); // DPI call to create transactor (called at
                                     // elaboration time as initialiser)

        bit report_available;

        // Function for getting a message from QUESTA_MVC. Returns 1 if a message was returned, 0 otherwise.
        import "DPI-C" questa_mvc_sv_get_report =  function bit get_report( input longint iface_ref,input longint recipient,
                                     output string category,     output string objectName,
                                     output string instanceName, output string error_no,
                                     output string typ,          output string mess );
        questa_mvc_reporter endPoint[longint];
        initial report_available = 0;

        always @report_available
        begin
            longint recipient;
            string category;
            string objectName;
            string instanceName;
            string severity;
            string mess;
            string error_no;

            if ( endPoint.first( recipient ) )
              begin
                do
                  begin
                      while ( get_report( _interface_ref, recipient, category, objectName, instanceName, error_no, severity, mess ) )
                        begin
                          endPoint[recipient].report_message( category, "axi", 0, objectName, instanceName, error_no, severity, mess );
                        end
                  end
                while (endPoint.next(recipient));
              end
            report_available = 0;
        end

        import "DPI-C" context questa_mvc_register_end_point = function void questa_mvc_register_end_point( input longint iface_ref, input longint as_end, input string name );

        // A function for registering a reporter to capture any reports coming from as_end
        function automatic void register_end_point( input longint as_end, input questa_mvc_reporter rep = null );
            if ( rep != null )
              begin
                if ( ( rep.name == "" ) || ( rep.name == "NULL" ) )
                  begin
                    $display("Error: %m: Reporter passed to register_end_point has a reserved name. Neither an empty string nor the string 'NULL' can be used.");
                  end
                else
                  begin
                    questa_mvc_register_end_point( _interface_ref, as_end, rep.name );
                    endPoint[as_end] = rep;
                  end
              end
            else
              begin
                questa_mvc_register_end_point( _interface_ref, as_end, "NULL" );
                endPoint.delete( as_end );
              end
        endfunction

    //-------------------------------------------------------------------------
    //
    // Group:- Registering Reports
    //
    //
    // The following methods are used to register a custom reporting object as
    // described in the MVC base library section, <Customizing Error-Reporting>.
    // 
    //-------------------------------------------------------------------------

    function void register_interface_reporter( input questa_mvc_reporter _rep = null );
        register_end_point( _interface_ref, _rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_master_reporter
    //
    // Function used to register a reporter for the <master> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the master end.
    //
    function void register_master_reporter
    (
        input questa_mvc_reporter rep = null
    );
        register_end_point( axi_master_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_slave_reporter
    //
    // Function used to register a reporter for the <slave> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the slave end.
    //
    function void register_slave_reporter
    (
        input questa_mvc_reporter rep = null
    );
        register_end_point( axi_slave_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_clock_source_reporter
    //
    // Function used to register a reporter for the <clock_source> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the clock_source end.
    //
    function void register_clock_source_reporter
    (
        input questa_mvc_reporter rep = null
    );
        register_end_point( axi_clock_source_end, rep );
    endfunction

    //-------------------------------------------------------------------------
    // Function:- register_reset_source_reporter
    //
    // Function used to register a reporter for the <reset_source> end of the
    // <axi> interface. See <Customizing Error-Reporting> for a
    // description of creating, customising and using reporters.
    //
    // Arguments:
    //    rep - The reporter to be used for the reset_source end.
    //
    function void register_reset_source_reporter
    (
        input questa_mvc_reporter rep = null
    );
        register_end_point( axi_reset_source_end, rep );
    endfunction


    //-------------------------------------------------------------------------
    //
    // Group:- BFM Utility/Convenience Methods
    //
    // This is the group of utility functions provided by the QVIP BFM to
    // communicate from the SV world to the QVIP BFM.
    // This set of APIs can be used to either get status/statistics
    // information from the BFM or to set values in a particular database 
    // in the BFM. Please refer to individual functions for more information.
    //
    //-------------------------------------------------------------------------

    export "DPI-C" axi_get_temp_static_fn_rd_txn_valid_lanes_valid_lanes = function axi_get_temp_static_fn_rd_txn_valid_lanes_valid_lanes;
    export "DPI-C" axi_set_temp_static_fn_rd_txn_valid_lanes_valid_lanes = function axi_set_temp_static_fn_rd_txn_valid_lanes_valid_lanes;
    bit [((AXI_RDATA_WIDTH / 8) - 1):0] temp_static_fn_rd_txn_valid_lanes_valid_lanes [];
    function void axi_get_temp_static_fn_rd_txn_valid_lanes_valid_lanes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_fn_rd_txn_valid_lanes_valid_lanes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_fn_rd_txn_valid_lanes_valid_lanes( input int _d1, input int _d2, input bit _value );
        temp_static_fn_rd_txn_valid_lanes_valid_lanes[_d1][_d2] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_rd_txn_valid_lanes
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get valid strobes/lanes value for each of the read data beat
    //     at end of read transaction.
    // 
    //     Please note that this function should be called after completion of a read
    //     transaction.
    // 
    //     Output of the function:
    //     valid_lanes - Valid strobes value for each read data beat
    //    
    function automatic void fn_rd_txn_valid_lanes
    (
        ref bit [((AXI_RDATA_WIDTH / 8) - 1):0] valid_lanes []
    );
        temp_static_fn_rd_txn_valid_lanes_valid_lanes = new[valid_lanes.size()];
         fn_rd_txn_valid_lanes_C();
        valid_lanes = temp_static_fn_rd_txn_valid_lanes_valid_lanes;
    endfunction

    export "DPI-C" axi_get_temp_static_fn_get_wdata_phase_info_id = function axi_get_temp_static_fn_get_wdata_phase_info_id;
    export "DPI-C" axi_set_temp_static_fn_get_wdata_phase_info_id = function axi_set_temp_static_fn_get_wdata_phase_info_id;
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_fn_get_wdata_phase_info_id;
    function void axi_get_temp_static_fn_get_wdata_phase_info_id( input int _d1, output bit  _value );
        _value = temp_static_fn_get_wdata_phase_info_id[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_wdata_phase_info_id( input int _d1, input bit  _value );
        temp_static_fn_get_wdata_phase_info_id[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_get_wdata_phase_info_beat_addr = function axi_get_temp_static_fn_get_wdata_phase_info_beat_addr;
    export "DPI-C" axi_set_temp_static_fn_get_wdata_phase_info_beat_addr = function axi_set_temp_static_fn_get_wdata_phase_info_beat_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_get_wdata_phase_info_beat_addr;
    function void axi_get_temp_static_fn_get_wdata_phase_info_beat_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_get_wdata_phase_info_beat_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_wdata_phase_info_beat_addr( input int _d1, input bit  _value );
        temp_static_fn_get_wdata_phase_info_beat_addr[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_get_wdata_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get information corresponding to a write data beat.
    // 
    //     Input:
    //     id         - ID of the write data beat
    //     wdata_last - assigned to ~last~ attribute of the write data beat
    // 
    //     Output:
    //     waddr_rcvd   - Indicates if corresponding write address phase is received
    //     burst_length - Burst length attribute of the corresponding address phase
    //     beat_num     - Write data beat number of the corresponding write data burst
    //     beat_addr    - Corresponding beat address
    // 
    //     Please note that this function should be called at the completion of write
    //     data beat.
    //    
    function automatic void fn_get_wdata_phase_info
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit wdata_last,
        inout bit waddr_rcvd,
        output bit [3:0] burst_length,
        output int beat_num,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  beat_addr
    );
        temp_static_fn_get_wdata_phase_info_id = id;
         fn_get_wdata_phase_info_C(wdata_last,waddr_rcvd,burst_length,beat_num);
        beat_addr = temp_static_fn_get_wdata_phase_info_beat_addr;
    endfunction

    export "DPI-C" axi_get_temp_static_fn_get_wresp_phase_info_wresp_corr_addr = function axi_get_temp_static_fn_get_wresp_phase_info_wresp_corr_addr;
    export "DPI-C" axi_set_temp_static_fn_get_wresp_phase_info_wresp_corr_addr = function axi_set_temp_static_fn_get_wresp_phase_info_wresp_corr_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_get_wresp_phase_info_wresp_corr_addr;
    function void axi_get_temp_static_fn_get_wresp_phase_info_wresp_corr_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_get_wresp_phase_info_wresp_corr_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_wresp_phase_info_wresp_corr_addr( input int _d1, input bit  _value );
        temp_static_fn_get_wresp_phase_info_wresp_corr_addr[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_get_wresp_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get address attribute of write address phase corresponding
    //     to write response phase that just completed.
    // 
    //     Please note that this function should be called after completion of a write
    //     response phase.
    // 
    //     Output of the function:
    //     wresp_corr_addr - ~addr~ attribute of the address phase corresponding to
    //                       this write response phase
    //    
    function automatic void fn_get_wresp_phase_info
    (
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  wresp_corr_addr
    );
         fn_get_wresp_phase_info_C();
        wresp_corr_addr = temp_static_fn_get_wresp_phase_info_wresp_corr_addr;
    endfunction

    export "DPI-C" axi_get_temp_static_fn_get_rdata_phase_info_id = function axi_get_temp_static_fn_get_rdata_phase_info_id;
    export "DPI-C" axi_set_temp_static_fn_get_rdata_phase_info_id = function axi_set_temp_static_fn_get_rdata_phase_info_id;
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_fn_get_rdata_phase_info_id;
    function void axi_get_temp_static_fn_get_rdata_phase_info_id( input int _d1, output bit  _value );
        _value = temp_static_fn_get_rdata_phase_info_id[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_rdata_phase_info_id( input int _d1, input bit  _value );
        temp_static_fn_get_rdata_phase_info_id[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_get_rdata_phase_info_beat_strobes = function axi_get_temp_static_fn_get_rdata_phase_info_beat_strobes;
    export "DPI-C" axi_set_temp_static_fn_get_rdata_phase_info_beat_strobes = function axi_set_temp_static_fn_get_rdata_phase_info_beat_strobes;
    bit [((AXI_RDATA_WIDTH / 8) - 1):0]  temp_static_fn_get_rdata_phase_info_beat_strobes;
    function void axi_get_temp_static_fn_get_rdata_phase_info_beat_strobes( input int _d1, output bit  _value );
        _value = temp_static_fn_get_rdata_phase_info_beat_strobes[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_rdata_phase_info_beat_strobes( input int _d1, input bit  _value );
        temp_static_fn_get_rdata_phase_info_beat_strobes[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_get_rdata_phase_info_beat_addr = function axi_get_temp_static_fn_get_rdata_phase_info_beat_addr;
    export "DPI-C" axi_set_temp_static_fn_get_rdata_phase_info_beat_addr = function axi_set_temp_static_fn_get_rdata_phase_info_beat_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_get_rdata_phase_info_beat_addr;
    function void axi_get_temp_static_fn_get_rdata_phase_info_beat_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_get_rdata_phase_info_beat_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_rdata_phase_info_beat_addr( input int _d1, input bit  _value );
        temp_static_fn_get_rdata_phase_info_beat_addr[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_get_rdata_phase_info_txn_addr = function axi_get_temp_static_fn_get_rdata_phase_info_txn_addr;
    export "DPI-C" axi_set_temp_static_fn_get_rdata_phase_info_txn_addr = function axi_set_temp_static_fn_get_rdata_phase_info_txn_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_get_rdata_phase_info_txn_addr;
    function void axi_get_temp_static_fn_get_rdata_phase_info_txn_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_get_rdata_phase_info_txn_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_get_rdata_phase_info_txn_addr( input int _d1, input bit  _value );
        temp_static_fn_get_rdata_phase_info_txn_addr[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_get_rdata_phase_info
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    //     A function to get information corresponding to a read data beat.
    // 
    //     Input:
    //     id         - ID of the read data beat
    // 
    //     Output:
    //     burst_length - Burst length attribute of the corresponding read address phase
    //     beat_num     - Read data beat number of the corresponding read data burst
    //     beat_strobes - Valid lanes in the read data beat
    //     beat_addr    - Corresponding beat address
    // 
    //     Please note that this function should be called at the completion of read
    //     data beat.
    //    
    function automatic void fn_get_rdata_phase_info
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit rdata_last,
        output bit [3:0] burst_length,
        output int beat_num,
        output bit [((AXI_RDATA_WIDTH / 8) - 1):0]  beat_strobes,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  beat_addr,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  txn_addr
    );
        temp_static_fn_get_rdata_phase_info_id = id;
         fn_get_rdata_phase_info_C(rdata_last,burst_length,beat_num);
        beat_strobes = temp_static_fn_get_rdata_phase_info_beat_strobes;
        beat_addr = temp_static_fn_get_rdata_phase_info_beat_addr;
        txn_addr = temp_static_fn_get_rdata_phase_info_txn_addr;
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_get_max_os_per_id
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function gets the maximum number of outstanding write phases of a particular ID
    // from among all AWID, WID values.
    //  
    // Inputs:
    // max_waddr_os - The maximum number of address phases outstanding from among all AWID
    // max_wdata_os - The maximum number of data bursts outstanding from among all WID
    // 
    // For example, 5 write address phases are outstanding with ID 3, and 
    // 7 write address phases are outstanding with ID 2. No other address phase is there
    // and 0 write data phases are received.
    // 
    // The return values would be such that:
    // max_waddr_os = 7
    // max_wdata_os = 0
    // 
    function automatic void fn_get_max_os_per_id
    (
        output int max_waddr_os,
        output int max_wdata_os
    );
         fn_get_max_os_per_id_C(max_waddr_os,max_wdata_os);
    endfunction

    export "DPI-C" axi_get_temp_static_get_rw_txns_in_prog_id = function axi_get_temp_static_get_rw_txns_in_prog_id;
    export "DPI-C" axi_set_temp_static_get_rw_txns_in_prog_id = function axi_set_temp_static_get_rw_txns_in_prog_id;
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_get_rw_txns_in_prog_id;
    function void axi_get_temp_static_get_rw_txns_in_prog_id( input int _d1, output bit  _value );
        _value = temp_static_get_rw_txns_in_prog_id[_d1];
    endfunction
    function void axi_set_temp_static_get_rw_txns_in_prog_id( input int _d1, input bit  _value );
        temp_static_get_rw_txns_in_prog_id[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: get_rw_txns_in_prog
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function gets the number of various outstanding transactions at a time.
    // 
    // Inputs:
    // id  - The AWID/ARID/WID of the transaction whose details are required.
    // txn_counts - The statistics of the number of outstanding transactions
    function automatic void get_rw_txns_in_prog
    (
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_rw_txn_counts_s txn_counts
    );
        temp_static_get_rw_txns_in_prog_id = id;
         get_rw_txns_in_prog_C(txn_counts);
    endfunction

    export "DPI-C" axi_get_temp_static_fn_add_addr_map_entry_addr = function axi_get_temp_static_fn_add_addr_map_entry_addr;
    export "DPI-C" axi_set_temp_static_fn_add_addr_map_entry_addr = function axi_set_temp_static_fn_add_addr_map_entry_addr;
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_fn_add_addr_map_entry_addr;
    function void axi_get_temp_static_fn_add_addr_map_entry_addr( input int _d1, output bit  _value );
        _value = temp_static_fn_add_addr_map_entry_addr[_d1];
    endfunction
    function void axi_set_temp_static_fn_add_addr_map_entry_addr( input int _d1, input bit  _value );
        temp_static_fn_add_addr_map_entry_addr[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_add_addr_map_entry
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets address map fields inside internal BFM. 
    // 
    // Inputs:
    // region - Region name 
    // addr - Start address of region
    // size - Size of address region
    function automatic void fn_add_addr_map_entry
    (
        input string region,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input longint unsigned size
    );
        temp_static_fn_add_addr_map_entry_addr = addr;
         fn_add_addr_map_entry_C(region,size);
    endfunction

    export "DPI-C" axi_get_temp_static_fn_add_wr_delay_data2data = function axi_get_temp_static_fn_add_wr_delay_data2data;
    export "DPI-C" axi_set_temp_static_fn_add_wr_delay_data2data = function axi_set_temp_static_fn_add_wr_delay_data2data;
    int unsigned temp_static_fn_add_wr_delay_data2data[];
    function void axi_get_temp_static_fn_add_wr_delay_data2data( input int _d1, output int unsigned _value );
        _value = temp_static_fn_add_wr_delay_data2data[_d1];
    endfunction
    function void axi_set_temp_static_fn_add_wr_delay_data2data( input int _d1, input int unsigned _value );
        temp_static_fn_add_wr_delay_data2data[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_add_wr_delay
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets delay values for write address-data pair and 
    // between write data beats, initiated by master end. 
    // 
    // Inputs:
    // region - Region value for which write delays are to be inserted
    // id - Write transaction's id (AWID) for which delays are to be inserted
    // addr2data - Delays to be inserted between write address and data phase.
    // data2data - Delays to be inserted between data beats
    function automatic void fn_add_wr_delay
    (
        input string region,
        input bit [17:0] id,
        input int unsigned addr2data,
        ref int unsigned data2data[]
    );
        int tmp_data2data_DIMS0;
        tmp_data2data_DIMS0 = data2data.size();
        temp_static_fn_add_wr_delay_data2data = data2data;
         fn_add_wr_delay_C(region,id,addr2data,tmp_data2data_DIMS0);
    endfunction

    //-------------------------------------------------------------------------
    // Function: fn_delete_wr_delay
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function deletes delay values for a region-id pair
    // 
    // Inputs:
    // region - Region value for which write delays are to be inserted
    // id - Write transaction's id (AWID) for which delays are to be inserted
    // addr2data - Delays to be inserted between write address and data phase.
    // data2data - Delays to be inserted between data beats
    function automatic void fn_delete_wr_delay
    (
        input string region,
        input bit [17:0] id
    );
         fn_delete_wr_delay_C(region,id);
    endfunction

    export "DPI-C" axi_get_temp_static_fn_set_wr_def_delays_min_data2data = function axi_get_temp_static_fn_set_wr_def_delays_min_data2data;
    export "DPI-C" axi_set_temp_static_fn_set_wr_def_delays_min_data2data = function axi_set_temp_static_fn_set_wr_def_delays_min_data2data;
    int unsigned temp_static_fn_set_wr_def_delays_min_data2data[];
    function void axi_get_temp_static_fn_set_wr_def_delays_min_data2data( input int _d1, output int unsigned _value );
        _value = temp_static_fn_set_wr_def_delays_min_data2data[_d1];
    endfunction
    function void axi_set_temp_static_fn_set_wr_def_delays_min_data2data( input int _d1, input int unsigned _value );
        temp_static_fn_set_wr_def_delays_min_data2data[_d1] = _value;
    endfunction
    export "DPI-C" axi_get_temp_static_fn_set_wr_def_delays_max_data2data = function axi_get_temp_static_fn_set_wr_def_delays_max_data2data;
    export "DPI-C" axi_set_temp_static_fn_set_wr_def_delays_max_data2data = function axi_set_temp_static_fn_set_wr_def_delays_max_data2data;
    int unsigned temp_static_fn_set_wr_def_delays_max_data2data[];
    function void axi_get_temp_static_fn_set_wr_def_delays_max_data2data( input int _d1, output int unsigned _value );
        _value = temp_static_fn_set_wr_def_delays_max_data2data[_d1];
    endfunction
    function void axi_set_temp_static_fn_set_wr_def_delays_max_data2data( input int _d1, input int unsigned _value );
        temp_static_fn_set_wr_def_delays_max_data2data[_d1] = _value;
    endfunction
    //-------------------------------------------------------------------------
    // Function: fn_set_wr_def_delays
    //-------------------------------------------------------------------------
    // ---------------------------------------------------------------------------
    // This function sets default delay values for write address-data pair and data beats 
    // initiated by master end between input max. and min. values. In case non-randomized 
    // default value is desired, user can set max. and min. to same value.
    // 
    // Inputs:
    // min_addr2data - Minimum value of default delays to be inserted between write address and data phase.
    // min_data2data - Minimum value of default delays to be inserted between data beats
    // max_addr2data - Maximum value of default delays to be inserted between write address and data phase.
    // max_data2data - Maximum value of default delays to be inserted between data beats
    function automatic void fn_set_wr_def_delays
    (
        input int unsigned min_addr2data,
        ref int unsigned min_data2data[],
        input int unsigned max_addr2data,
        ref int unsigned max_data2data[]
    );
        int tmp_min_data2data_DIMS0;
        int tmp_max_data2data_DIMS0;
        tmp_min_data2data_DIMS0 = min_data2data.size();
        tmp_max_data2data_DIMS0 = max_data2data.size();
        temp_static_fn_set_wr_def_delays_min_data2data = min_data2data;
        temp_static_fn_set_wr_def_delays_max_data2data = max_data2data;
         fn_set_wr_def_delays_C(min_addr2data,tmp_min_data2data_DIMS0,max_addr2data,tmp_max_data2data_DIMS0);
    endfunction

    // Declare user visible wires variables, for non-continuous assignments.
    logic m_ACLK = 'z;
    logic m_ARESETn = 'z;
    logic m_AWVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  m_AWADDR = 'z;
    logic [3:0] m_AWLEN = 'z;
    logic [2:0] m_AWSIZE = 'z;
    logic [1:0] m_AWBURST = 'z;
    logic [1:0] m_AWLOCK = 'z;
    logic [3:0] m_AWCACHE = 'z;
    logic [2:0] m_AWPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_AWID = 'z;
    logic m_AWREADY = 'z;
    logic [7:0] m_AWUSER = 'z;
    logic m_ARVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  m_ARADDR = 'z;
    logic [3:0] m_ARLEN = 'z;
    logic [2:0] m_ARSIZE = 'z;
    logic [1:0] m_ARBURST = 'z;
    logic [1:0] m_ARLOCK = 'z;
    logic [3:0] m_ARCACHE = 'z;
    logic [2:0] m_ARPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_ARID = 'z;
    logic m_ARREADY = 'z;
    logic [7:0] m_ARUSER = 'z;
    logic m_RVALID = 'z;
    logic m_RLAST = 'z;
    logic [((AXI_RDATA_WIDTH) - 1):0]  m_RDATA = 'z;
    logic [1:0] m_RRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_RID = 'z;
    logic m_RREADY = 'z;
    logic [7:0] m_RUSER = 'z;
    logic m_WVALID = 'z;
    logic m_WLAST = 'z;
    logic [((AXI_WDATA_WIDTH) - 1):0]  m_WDATA = 'z;
    logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  m_WSTRB = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_WID = 'z;
    logic m_WREADY = 'z;
    logic [7:0] m_WUSER = 'z;
    logic m_BVALID = 'z;
    logic [1:0] m_BRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  m_BID = 'z;
    logic m_BREADY = 'z;
    logic [7:0] m_BUSER = 'z;

    // Forces a sweep through the wire change checkers at time 0 to get around
    // process kick-off order unknowns
    bit _check_t0_values;
    always_comb _check_t0_values = 1;

    // handle control
    longint last_handle = 0;

    longint last_start_time = 0;

    longint last_end_time = 0;

    export "DPI-C" axi_set_last_handle_and_times = function set_last_handle_and_times;

    function void set_last_handle_and_times(longint _handle, longint _start, longint _end);
        last_handle = _handle;
        last_start_time = _start;
        last_end_time = _end;
    endfunction


    function longint get_last_handle();
        return last_handle;
    endfunction


    function longint get_last_start_time();
        return last_start_time;
    endfunction


    function longint get_last_end_time();
        return last_end_time;
    endfunction


    //-------------------------------------------------------------------------
    // Tasks to wait for a number of specified edges on a wire
    //-------------------------------------------------------------------------


    //------------------------------------------------------------------------------
    // Function:- wait_for_ACLK
    //     Wait for the specified change on wire <axi::ACLK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ACLK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ACLK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ACLK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ACLK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ACLK === 0 );
                    @( ACLK );
                end
                while ( ACLK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ACLK === 1 );
                    @( ACLK );
                end
                while ( ACLK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARESETn
    //     Wait for the specified change on wire <axi::ARESETn>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARESETn( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARESETn);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARESETn);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARESETn);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARESETn === 0 );
                    @( ARESETn );
                end
                while ( ARESETn !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARESETn === 1 );
                    @( ARESETn );
                end
                while ( ARESETn !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWVALID
    //     Wait for the specified change on wire <axi::AWVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWVALID === 0 );
                    @( AWVALID );
                end
                while ( AWVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWVALID === 1 );
                    @( AWVALID );
                end
                while ( AWVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWADDR
    //     Wait for the specified change on wire <axi::AWADDR>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWADDR( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWADDR);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWADDR);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWADDR);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWADDR === 0 );
                    @( AWADDR );
                end
                while ( AWADDR !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWADDR === 1 );
                    @( AWADDR );
                end
                while ( AWADDR !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWADDR_index1
    //     Wait for the specified change on wire <axi::AWADDR>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWADDR_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWADDR[_this_dot_1] === 0 );
                    @( AWADDR[_this_dot_1] );
                end
                while ( AWADDR[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWADDR[_this_dot_1] === 1 );
                    @( AWADDR[_this_dot_1] );
                end
                while ( AWADDR[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLEN
    //     Wait for the specified change on wire <axi::AWLEN>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLEN( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLEN);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLEN);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLEN);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLEN === 0 );
                    @( AWLEN );
                end
                while ( AWLEN !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLEN === 1 );
                    @( AWLEN );
                end
                while ( AWLEN !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLEN_index1
    //     Wait for the specified change on wire <axi::AWLEN>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLEN_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLEN[_this_dot_1] === 0 );
                    @( AWLEN[_this_dot_1] );
                end
                while ( AWLEN[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLEN[_this_dot_1] === 1 );
                    @( AWLEN[_this_dot_1] );
                end
                while ( AWLEN[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWSIZE
    //     Wait for the specified change on wire <axi::AWSIZE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWSIZE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWSIZE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWSIZE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWSIZE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWSIZE === 0 );
                    @( AWSIZE );
                end
                while ( AWSIZE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWSIZE === 1 );
                    @( AWSIZE );
                end
                while ( AWSIZE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWSIZE_index1
    //     Wait for the specified change on wire <axi::AWSIZE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWSIZE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWSIZE[_this_dot_1] === 0 );
                    @( AWSIZE[_this_dot_1] );
                end
                while ( AWSIZE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWSIZE[_this_dot_1] === 1 );
                    @( AWSIZE[_this_dot_1] );
                end
                while ( AWSIZE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWBURST
    //     Wait for the specified change on wire <axi::AWBURST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWBURST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWBURST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWBURST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWBURST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWBURST === 0 );
                    @( AWBURST );
                end
                while ( AWBURST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWBURST === 1 );
                    @( AWBURST );
                end
                while ( AWBURST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWBURST_index1
    //     Wait for the specified change on wire <axi::AWBURST>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWBURST_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWBURST[_this_dot_1] === 0 );
                    @( AWBURST[_this_dot_1] );
                end
                while ( AWBURST[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWBURST[_this_dot_1] === 1 );
                    @( AWBURST[_this_dot_1] );
                end
                while ( AWBURST[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLOCK
    //     Wait for the specified change on wire <axi::AWLOCK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLOCK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLOCK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLOCK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLOCK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLOCK === 0 );
                    @( AWLOCK );
                end
                while ( AWLOCK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLOCK === 1 );
                    @( AWLOCK );
                end
                while ( AWLOCK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWLOCK_index1
    //     Wait for the specified change on wire <axi::AWLOCK>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWLOCK_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWLOCK[_this_dot_1] === 0 );
                    @( AWLOCK[_this_dot_1] );
                end
                while ( AWLOCK[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWLOCK[_this_dot_1] === 1 );
                    @( AWLOCK[_this_dot_1] );
                end
                while ( AWLOCK[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWCACHE
    //     Wait for the specified change on wire <axi::AWCACHE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWCACHE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWCACHE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWCACHE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWCACHE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWCACHE === 0 );
                    @( AWCACHE );
                end
                while ( AWCACHE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWCACHE === 1 );
                    @( AWCACHE );
                end
                while ( AWCACHE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWCACHE_index1
    //     Wait for the specified change on wire <axi::AWCACHE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWCACHE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWCACHE[_this_dot_1] === 0 );
                    @( AWCACHE[_this_dot_1] );
                end
                while ( AWCACHE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWCACHE[_this_dot_1] === 1 );
                    @( AWCACHE[_this_dot_1] );
                end
                while ( AWCACHE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWPROT
    //     Wait for the specified change on wire <axi::AWPROT>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWPROT( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWPROT);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWPROT);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWPROT);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWPROT === 0 );
                    @( AWPROT );
                end
                while ( AWPROT !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWPROT === 1 );
                    @( AWPROT );
                end
                while ( AWPROT !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWPROT_index1
    //     Wait for the specified change on wire <axi::AWPROT>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWPROT_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWPROT[_this_dot_1] === 0 );
                    @( AWPROT[_this_dot_1] );
                end
                while ( AWPROT[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWPROT[_this_dot_1] === 1 );
                    @( AWPROT[_this_dot_1] );
                end
                while ( AWPROT[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWID
    //     Wait for the specified change on wire <axi::AWID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWID === 0 );
                    @( AWID );
                end
                while ( AWID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWID === 1 );
                    @( AWID );
                end
                while ( AWID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWID_index1
    //     Wait for the specified change on wire <axi::AWID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWID[_this_dot_1] === 0 );
                    @( AWID[_this_dot_1] );
                end
                while ( AWID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWID[_this_dot_1] === 1 );
                    @( AWID[_this_dot_1] );
                end
                while ( AWID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWREADY
    //     Wait for the specified change on wire <axi::AWREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWREADY === 0 );
                    @( AWREADY );
                end
                while ( AWREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWREADY === 1 );
                    @( AWREADY );
                end
                while ( AWREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWUSER
    //     Wait for the specified change on wire <axi::AWUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWUSER === 0 );
                    @( AWUSER );
                end
                while ( AWUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWUSER === 1 );
                    @( AWUSER );
                end
                while ( AWUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_AWUSER_index1
    //     Wait for the specified change on wire <axi::AWUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_AWUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        AWUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( AWUSER[_this_dot_1] === 0 );
                    @( AWUSER[_this_dot_1] );
                end
                while ( AWUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( AWUSER[_this_dot_1] === 1 );
                    @( AWUSER[_this_dot_1] );
                end
                while ( AWUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARVALID
    //     Wait for the specified change on wire <axi::ARVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARVALID === 0 );
                    @( ARVALID );
                end
                while ( ARVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARVALID === 1 );
                    @( ARVALID );
                end
                while ( ARVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARADDR
    //     Wait for the specified change on wire <axi::ARADDR>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARADDR( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARADDR);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARADDR);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARADDR);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARADDR === 0 );
                    @( ARADDR );
                end
                while ( ARADDR !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARADDR === 1 );
                    @( ARADDR );
                end
                while ( ARADDR !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARADDR_index1
    //     Wait for the specified change on wire <axi::ARADDR>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARADDR_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARADDR[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARADDR[_this_dot_1] === 0 );
                    @( ARADDR[_this_dot_1] );
                end
                while ( ARADDR[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARADDR[_this_dot_1] === 1 );
                    @( ARADDR[_this_dot_1] );
                end
                while ( ARADDR[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLEN
    //     Wait for the specified change on wire <axi::ARLEN>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLEN( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLEN);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLEN);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLEN);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLEN === 0 );
                    @( ARLEN );
                end
                while ( ARLEN !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLEN === 1 );
                    @( ARLEN );
                end
                while ( ARLEN !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLEN_index1
    //     Wait for the specified change on wire <axi::ARLEN>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLEN_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLEN[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLEN[_this_dot_1] === 0 );
                    @( ARLEN[_this_dot_1] );
                end
                while ( ARLEN[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLEN[_this_dot_1] === 1 );
                    @( ARLEN[_this_dot_1] );
                end
                while ( ARLEN[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARSIZE
    //     Wait for the specified change on wire <axi::ARSIZE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARSIZE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARSIZE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARSIZE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARSIZE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARSIZE === 0 );
                    @( ARSIZE );
                end
                while ( ARSIZE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARSIZE === 1 );
                    @( ARSIZE );
                end
                while ( ARSIZE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARSIZE_index1
    //     Wait for the specified change on wire <axi::ARSIZE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARSIZE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARSIZE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARSIZE[_this_dot_1] === 0 );
                    @( ARSIZE[_this_dot_1] );
                end
                while ( ARSIZE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARSIZE[_this_dot_1] === 1 );
                    @( ARSIZE[_this_dot_1] );
                end
                while ( ARSIZE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARBURST
    //     Wait for the specified change on wire <axi::ARBURST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARBURST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARBURST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARBURST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARBURST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARBURST === 0 );
                    @( ARBURST );
                end
                while ( ARBURST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARBURST === 1 );
                    @( ARBURST );
                end
                while ( ARBURST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARBURST_index1
    //     Wait for the specified change on wire <axi::ARBURST>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARBURST_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARBURST[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARBURST[_this_dot_1] === 0 );
                    @( ARBURST[_this_dot_1] );
                end
                while ( ARBURST[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARBURST[_this_dot_1] === 1 );
                    @( ARBURST[_this_dot_1] );
                end
                while ( ARBURST[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLOCK
    //     Wait for the specified change on wire <axi::ARLOCK>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLOCK( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLOCK);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLOCK);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLOCK);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLOCK === 0 );
                    @( ARLOCK );
                end
                while ( ARLOCK !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLOCK === 1 );
                    @( ARLOCK );
                end
                while ( ARLOCK !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARLOCK_index1
    //     Wait for the specified change on wire <axi::ARLOCK>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARLOCK_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARLOCK[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARLOCK[_this_dot_1] === 0 );
                    @( ARLOCK[_this_dot_1] );
                end
                while ( ARLOCK[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARLOCK[_this_dot_1] === 1 );
                    @( ARLOCK[_this_dot_1] );
                end
                while ( ARLOCK[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARCACHE
    //     Wait for the specified change on wire <axi::ARCACHE>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARCACHE( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARCACHE);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARCACHE);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARCACHE);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARCACHE === 0 );
                    @( ARCACHE );
                end
                while ( ARCACHE !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARCACHE === 1 );
                    @( ARCACHE );
                end
                while ( ARCACHE !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARCACHE_index1
    //     Wait for the specified change on wire <axi::ARCACHE>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARCACHE_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARCACHE[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARCACHE[_this_dot_1] === 0 );
                    @( ARCACHE[_this_dot_1] );
                end
                while ( ARCACHE[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARCACHE[_this_dot_1] === 1 );
                    @( ARCACHE[_this_dot_1] );
                end
                while ( ARCACHE[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARPROT
    //     Wait for the specified change on wire <axi::ARPROT>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARPROT( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARPROT);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARPROT);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARPROT);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARPROT === 0 );
                    @( ARPROT );
                end
                while ( ARPROT !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARPROT === 1 );
                    @( ARPROT );
                end
                while ( ARPROT !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARPROT_index1
    //     Wait for the specified change on wire <axi::ARPROT>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARPROT_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARPROT[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARPROT[_this_dot_1] === 0 );
                    @( ARPROT[_this_dot_1] );
                end
                while ( ARPROT[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARPROT[_this_dot_1] === 1 );
                    @( ARPROT[_this_dot_1] );
                end
                while ( ARPROT[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARID
    //     Wait for the specified change on wire <axi::ARID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARID === 0 );
                    @( ARID );
                end
                while ( ARID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARID === 1 );
                    @( ARID );
                end
                while ( ARID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARID_index1
    //     Wait for the specified change on wire <axi::ARID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARID[_this_dot_1] === 0 );
                    @( ARID[_this_dot_1] );
                end
                while ( ARID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARID[_this_dot_1] === 1 );
                    @( ARID[_this_dot_1] );
                end
                while ( ARID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARREADY
    //     Wait for the specified change on wire <axi::ARREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARREADY === 0 );
                    @( ARREADY );
                end
                while ( ARREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARREADY === 1 );
                    @( ARREADY );
                end
                while ( ARREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARUSER
    //     Wait for the specified change on wire <axi::ARUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARUSER === 0 );
                    @( ARUSER );
                end
                while ( ARUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARUSER === 1 );
                    @( ARUSER );
                end
                while ( ARUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_ARUSER_index1
    //     Wait for the specified change on wire <axi::ARUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_ARUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        ARUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( ARUSER[_this_dot_1] === 0 );
                    @( ARUSER[_this_dot_1] );
                end
                while ( ARUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( ARUSER[_this_dot_1] === 1 );
                    @( ARUSER[_this_dot_1] );
                end
                while ( ARUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RVALID
    //     Wait for the specified change on wire <axi::RVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RVALID === 0 );
                    @( RVALID );
                end
                while ( RVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RVALID === 1 );
                    @( RVALID );
                end
                while ( RVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RLAST
    //     Wait for the specified change on wire <axi::RLAST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RLAST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RLAST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RLAST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RLAST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RLAST === 0 );
                    @( RLAST );
                end
                while ( RLAST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RLAST === 1 );
                    @( RLAST );
                end
                while ( RLAST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RDATA
    //     Wait for the specified change on wire <axi::RDATA>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RDATA( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RDATA);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RDATA);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RDATA);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RDATA === 0 );
                    @( RDATA );
                end
                while ( RDATA !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RDATA === 1 );
                    @( RDATA );
                end
                while ( RDATA !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RDATA_index1
    //     Wait for the specified change on wire <axi::RDATA>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RDATA_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RDATA[_this_dot_1] === 0 );
                    @( RDATA[_this_dot_1] );
                end
                while ( RDATA[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RDATA[_this_dot_1] === 1 );
                    @( RDATA[_this_dot_1] );
                end
                while ( RDATA[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RRESP
    //     Wait for the specified change on wire <axi::RRESP>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RRESP( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RRESP);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RRESP);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RRESP);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RRESP === 0 );
                    @( RRESP );
                end
                while ( RRESP !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RRESP === 1 );
                    @( RRESP );
                end
                while ( RRESP !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RRESP_index1
    //     Wait for the specified change on wire <axi::RRESP>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RRESP_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RRESP[_this_dot_1] === 0 );
                    @( RRESP[_this_dot_1] );
                end
                while ( RRESP[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RRESP[_this_dot_1] === 1 );
                    @( RRESP[_this_dot_1] );
                end
                while ( RRESP[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RID
    //     Wait for the specified change on wire <axi::RID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RID === 0 );
                    @( RID );
                end
                while ( RID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RID === 1 );
                    @( RID );
                end
                while ( RID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RID_index1
    //     Wait for the specified change on wire <axi::RID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RID[_this_dot_1] === 0 );
                    @( RID[_this_dot_1] );
                end
                while ( RID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RID[_this_dot_1] === 1 );
                    @( RID[_this_dot_1] );
                end
                while ( RID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RREADY
    //     Wait for the specified change on wire <axi::RREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RREADY === 0 );
                    @( RREADY );
                end
                while ( RREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RREADY === 1 );
                    @( RREADY );
                end
                while ( RREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RUSER
    //     Wait for the specified change on wire <axi::RUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RUSER === 0 );
                    @( RUSER );
                end
                while ( RUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RUSER === 1 );
                    @( RUSER );
                end
                while ( RUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_RUSER_index1
    //     Wait for the specified change on wire <axi::RUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_RUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        RUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( RUSER[_this_dot_1] === 0 );
                    @( RUSER[_this_dot_1] );
                end
                while ( RUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( RUSER[_this_dot_1] === 1 );
                    @( RUSER[_this_dot_1] );
                end
                while ( RUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WVALID
    //     Wait for the specified change on wire <axi::WVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WVALID === 0 );
                    @( WVALID );
                end
                while ( WVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WVALID === 1 );
                    @( WVALID );
                end
                while ( WVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WLAST
    //     Wait for the specified change on wire <axi::WLAST>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WLAST( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WLAST);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WLAST);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WLAST);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WLAST === 0 );
                    @( WLAST );
                end
                while ( WLAST !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WLAST === 1 );
                    @( WLAST );
                end
                while ( WLAST !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WDATA
    //     Wait for the specified change on wire <axi::WDATA>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WDATA( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WDATA);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WDATA);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WDATA);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WDATA === 0 );
                    @( WDATA );
                end
                while ( WDATA !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WDATA === 1 );
                    @( WDATA );
                end
                while ( WDATA !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WDATA_index1
    //     Wait for the specified change on wire <axi::WDATA>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WDATA_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WDATA[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WDATA[_this_dot_1] === 0 );
                    @( WDATA[_this_dot_1] );
                end
                while ( WDATA[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WDATA[_this_dot_1] === 1 );
                    @( WDATA[_this_dot_1] );
                end
                while ( WDATA[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WSTRB
    //     Wait for the specified change on wire <axi::WSTRB>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WSTRB( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WSTRB);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WSTRB);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WSTRB);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WSTRB === 0 );
                    @( WSTRB );
                end
                while ( WSTRB !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WSTRB === 1 );
                    @( WSTRB );
                end
                while ( WSTRB !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WSTRB_index1
    //     Wait for the specified change on wire <axi::WSTRB>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WSTRB_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WSTRB[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WSTRB[_this_dot_1] === 0 );
                    @( WSTRB[_this_dot_1] );
                end
                while ( WSTRB[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WSTRB[_this_dot_1] === 1 );
                    @( WSTRB[_this_dot_1] );
                end
                while ( WSTRB[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WID
    //     Wait for the specified change on wire <axi::WID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WID === 0 );
                    @( WID );
                end
                while ( WID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WID === 1 );
                    @( WID );
                end
                while ( WID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WID_index1
    //     Wait for the specified change on wire <axi::WID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WID[_this_dot_1] === 0 );
                    @( WID[_this_dot_1] );
                end
                while ( WID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WID[_this_dot_1] === 1 );
                    @( WID[_this_dot_1] );
                end
                while ( WID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WREADY
    //     Wait for the specified change on wire <axi::WREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WREADY === 0 );
                    @( WREADY );
                end
                while ( WREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WREADY === 1 );
                    @( WREADY );
                end
                while ( WREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WUSER
    //     Wait for the specified change on wire <axi::WUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WUSER === 0 );
                    @( WUSER );
                end
                while ( WUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WUSER === 1 );
                    @( WUSER );
                end
                while ( WUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_WUSER_index1
    //     Wait for the specified change on wire <axi::WUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_WUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        WUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( WUSER[_this_dot_1] === 0 );
                    @( WUSER[_this_dot_1] );
                end
                while ( WUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( WUSER[_this_dot_1] === 1 );
                    @( WUSER[_this_dot_1] );
                end
                while ( WUSER[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BVALID
    //     Wait for the specified change on wire <axi::BVALID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BVALID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BVALID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BVALID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BVALID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BVALID === 0 );
                    @( BVALID );
                end
                while ( BVALID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BVALID === 1 );
                    @( BVALID );
                end
                while ( BVALID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BRESP
    //     Wait for the specified change on wire <axi::BRESP>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BRESP( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BRESP);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BRESP);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BRESP);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BRESP === 0 );
                    @( BRESP );
                end
                while ( BRESP !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BRESP === 1 );
                    @( BRESP );
                end
                while ( BRESP !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BRESP_index1
    //     Wait for the specified change on wire <axi::BRESP>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BRESP_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BRESP[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BRESP[_this_dot_1] === 0 );
                    @( BRESP[_this_dot_1] );
                end
                while ( BRESP[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BRESP[_this_dot_1] === 1 );
                    @( BRESP[_this_dot_1] );
                end
                while ( BRESP[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BID
    //     Wait for the specified change on wire <axi::BID>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BID( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BID);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BID);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BID);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BID === 0 );
                    @( BID );
                end
                while ( BID !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BID === 1 );
                    @( BID );
                end
                while ( BID !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BID_index1
    //     Wait for the specified change on wire <axi::BID>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BID_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BID[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BID[_this_dot_1] === 0 );
                    @( BID[_this_dot_1] );
                end
                while ( BID[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BID[_this_dot_1] === 1 );
                    @( BID[_this_dot_1] );
                end
                while ( BID[_this_dot_1] !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BREADY
    //     Wait for the specified change on wire <axi::BREADY>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BREADY( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BREADY);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BREADY);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BREADY);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BREADY === 0 );
                    @( BREADY );
                end
                while ( BREADY !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BREADY === 1 );
                    @( BREADY );
                end
                while ( BREADY !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BUSER
    //     Wait for the specified change on wire <axi::BUSER>.
    //
    // Arguments:
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BUSER( input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BUSER);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BUSER);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BUSER);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BUSER === 0 );
                    @( BUSER );
                end
                while ( BUSER !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BUSER === 1 );
                    @( BUSER );
                end
                while ( BUSER !== 0 );
            end
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_BUSER_index1
    //     Wait for the specified change on wire <axi::BUSER>.
    //
    // Arguments:
    //    _this_dot_1 - The array index for dimension 1.
    //     which_edge - The type of edge to wait for, one of <questa_mvc_edge>.
    //     count - The number of edges to wait for.
    //
    task automatic wait_for_BUSER_index1( input int _this_dot_1, input questa_mvc_edge which_edge, input int count = 1 );
        int i;
        for ( i=0; i<count; i++ )
        begin
            if      ( which_edge == QUESTA_MVC_POSEDGE     ) @(posedge BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_NEGEDGE     ) @(negedge BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_ANYEDGE     ) @(        BUSER[_this_dot_1]);
            else if ( which_edge == QUESTA_MVC_0_TO_1_EDGE )
            begin
                do
                begin
                    wait( BUSER[_this_dot_1] === 0 );
                    @( BUSER[_this_dot_1] );
                end
                while ( BUSER[_this_dot_1] !== 1 );
            end
            else if ( which_edge == QUESTA_MVC_1_TO_0_EDGE )
            begin
                do
                begin
                    wait( BUSER[_this_dot_1] === 1 );
                    @( BUSER[_this_dot_1] );
                end
                while ( BUSER[_this_dot_1] !== 0 );
            end
        end
    endtask

    //-------------------------------------------------------------------------
    // Tasks/functions to set/get wires
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- set_ACLK
    //-------------------------------------------------------------------------
    //     Set the value of wire <ACLK>.
    //
    // Parameters:
    //     ACLK_param - The value to set onto wire <ACLK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ACLK( logic ACLK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ACLK = ACLK_param;
        else
            m_ACLK <= ACLK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ACLK
    //-------------------------------------------------------------------------
    //     Get the value of wire <ACLK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ACLK>.
    //
    function automatic logic get_ACLK(  );
        return ACLK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARESETn
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARESETn>.
    //
    // Parameters:
    //     ARESETn_param - The value to set onto wire <ARESETn>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARESETn( logic ARESETn_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARESETn = ARESETn_param;
        else
            m_ARESETn <= ARESETn_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARESETn
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARESETn>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARESETn>.
    //
    function automatic logic get_ARESETn(  );
        return ARESETn;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWVALID>.
    //
    // Parameters:
    //     AWVALID_param - The value to set onto wire <AWVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWVALID( logic AWVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWVALID = AWVALID_param;
        else
            m_AWVALID <= AWVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWVALID>.
    //
    function automatic logic get_AWVALID(  );
        return AWVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWADDR
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWADDR>.
    //
    // Parameters:
    //     AWADDR_param - The value to set onto wire <AWADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWADDR( logic [((AXI_ADDRESS_WIDTH) - 1):0]  AWADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWADDR = AWADDR_param;
        else
            m_AWADDR <= AWADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWADDR_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWADDR_param - The value to set onto wire <AWADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWADDR_index1( int _this_dot_1, logic  AWADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWADDR[_this_dot_1] = AWADDR_param;
        else
            m_AWADDR[_this_dot_1] <= AWADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWADDR
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWADDR>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWADDR>.
    //
    function automatic logic [((AXI_ADDRESS_WIDTH) - 1):0]   get_AWADDR(  );
        return AWADDR;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWADDR_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWADDR>.
    //
    function automatic logic   get_AWADDR_index1( int _this_dot_1 );
        return AWADDR[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWLEN
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWLEN>.
    //
    // Parameters:
    //     AWLEN_param - The value to set onto wire <AWLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLEN( logic [3:0] AWLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLEN = AWLEN_param;
        else
            m_AWLEN <= AWLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWLEN_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWLEN_param - The value to set onto wire <AWLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLEN_index1( int _this_dot_1, logic  AWLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLEN[_this_dot_1] = AWLEN_param;
        else
            m_AWLEN[_this_dot_1] <= AWLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWLEN
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWLEN>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWLEN>.
    //
    function automatic logic [3:0]  get_AWLEN(  );
        return AWLEN;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWLEN_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWLEN>.
    //
    function automatic logic   get_AWLEN_index1( int _this_dot_1 );
        return AWLEN[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWSIZE
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWSIZE>.
    //
    // Parameters:
    //     AWSIZE_param - The value to set onto wire <AWSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWSIZE( logic [2:0] AWSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWSIZE = AWSIZE_param;
        else
            m_AWSIZE <= AWSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWSIZE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWSIZE_param - The value to set onto wire <AWSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWSIZE_index1( int _this_dot_1, logic  AWSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWSIZE[_this_dot_1] = AWSIZE_param;
        else
            m_AWSIZE[_this_dot_1] <= AWSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWSIZE
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWSIZE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWSIZE>.
    //
    function automatic logic [2:0]  get_AWSIZE(  );
        return AWSIZE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWSIZE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWSIZE>.
    //
    function automatic logic   get_AWSIZE_index1( int _this_dot_1 );
        return AWSIZE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWBURST
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWBURST>.
    //
    // Parameters:
    //     AWBURST_param - The value to set onto wire <AWBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWBURST( logic [1:0] AWBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWBURST = AWBURST_param;
        else
            m_AWBURST <= AWBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWBURST_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWBURST_param - The value to set onto wire <AWBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWBURST_index1( int _this_dot_1, logic  AWBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWBURST[_this_dot_1] = AWBURST_param;
        else
            m_AWBURST[_this_dot_1] <= AWBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWBURST
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWBURST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWBURST>.
    //
    function automatic logic [1:0]  get_AWBURST(  );
        return AWBURST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWBURST_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWBURST>.
    //
    function automatic logic   get_AWBURST_index1( int _this_dot_1 );
        return AWBURST[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWLOCK
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWLOCK>.
    //
    // Parameters:
    //     AWLOCK_param - The value to set onto wire <AWLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLOCK( logic [1:0] AWLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLOCK = AWLOCK_param;
        else
            m_AWLOCK <= AWLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWLOCK_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWLOCK_param - The value to set onto wire <AWLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWLOCK_index1( int _this_dot_1, logic  AWLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWLOCK[_this_dot_1] = AWLOCK_param;
        else
            m_AWLOCK[_this_dot_1] <= AWLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWLOCK
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWLOCK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWLOCK>.
    //
    function automatic logic [1:0]  get_AWLOCK(  );
        return AWLOCK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWLOCK_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWLOCK>.
    //
    function automatic logic   get_AWLOCK_index1( int _this_dot_1 );
        return AWLOCK[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWCACHE
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWCACHE>.
    //
    // Parameters:
    //     AWCACHE_param - The value to set onto wire <AWCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWCACHE( logic [3:0] AWCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWCACHE = AWCACHE_param;
        else
            m_AWCACHE <= AWCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWCACHE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWCACHE_param - The value to set onto wire <AWCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWCACHE_index1( int _this_dot_1, logic  AWCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWCACHE[_this_dot_1] = AWCACHE_param;
        else
            m_AWCACHE[_this_dot_1] <= AWCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWCACHE
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWCACHE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWCACHE>.
    //
    function automatic logic [3:0]  get_AWCACHE(  );
        return AWCACHE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWCACHE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWCACHE>.
    //
    function automatic logic   get_AWCACHE_index1( int _this_dot_1 );
        return AWCACHE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWPROT
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWPROT>.
    //
    // Parameters:
    //     AWPROT_param - The value to set onto wire <AWPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWPROT( logic [2:0] AWPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWPROT = AWPROT_param;
        else
            m_AWPROT <= AWPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWPROT_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWPROT_param - The value to set onto wire <AWPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWPROT_index1( int _this_dot_1, logic  AWPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWPROT[_this_dot_1] = AWPROT_param;
        else
            m_AWPROT[_this_dot_1] <= AWPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWPROT
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWPROT>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWPROT>.
    //
    function automatic logic [2:0]  get_AWPROT(  );
        return AWPROT;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWPROT_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWPROT>.
    //
    function automatic logic   get_AWPROT_index1( int _this_dot_1 );
        return AWPROT[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWID
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWID>.
    //
    // Parameters:
    //     AWID_param - The value to set onto wire <AWID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWID( logic [((AXI_ID_WIDTH) - 1):0]  AWID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWID = AWID_param;
        else
            m_AWID <= AWID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWID_param - The value to set onto wire <AWID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWID_index1( int _this_dot_1, logic  AWID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWID[_this_dot_1] = AWID_param;
        else
            m_AWID[_this_dot_1] <= AWID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWID
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_AWID(  );
        return AWID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWID>.
    //
    function automatic logic   get_AWID_index1( int _this_dot_1 );
        return AWID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWREADY>.
    //
    // Parameters:
    //     AWREADY_param - The value to set onto wire <AWREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWREADY( logic AWREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWREADY = AWREADY_param;
        else
            m_AWREADY <= AWREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWREADY>.
    //
    function automatic logic get_AWREADY(  );
        return AWREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_AWUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <AWUSER>.
    //
    // Parameters:
    //     AWUSER_param - The value to set onto wire <AWUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWUSER( logic [7:0] AWUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWUSER = AWUSER_param;
        else
            m_AWUSER <= AWUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_AWUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <AWUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     AWUSER_param - The value to set onto wire <AWUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_AWUSER_index1( int _this_dot_1, logic  AWUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_AWUSER[_this_dot_1] = AWUSER_param;
        else
            m_AWUSER[_this_dot_1] <= AWUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_AWUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <AWUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <AWUSER>.
    //
    function automatic logic [7:0]  get_AWUSER(  );
        return AWUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_AWUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <AWUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <AWUSER>.
    //
    function automatic logic   get_AWUSER_index1( int _this_dot_1 );
        return AWUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARVALID>.
    //
    // Parameters:
    //     ARVALID_param - The value to set onto wire <ARVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARVALID( logic ARVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARVALID = ARVALID_param;
        else
            m_ARVALID <= ARVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARVALID>.
    //
    function automatic logic get_ARVALID(  );
        return ARVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARADDR
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARADDR>.
    //
    // Parameters:
    //     ARADDR_param - The value to set onto wire <ARADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARADDR( logic [((AXI_ADDRESS_WIDTH) - 1):0]  ARADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARADDR = ARADDR_param;
        else
            m_ARADDR <= ARADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARADDR_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARADDR_param - The value to set onto wire <ARADDR>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARADDR_index1( int _this_dot_1, logic  ARADDR_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARADDR[_this_dot_1] = ARADDR_param;
        else
            m_ARADDR[_this_dot_1] <= ARADDR_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARADDR
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARADDR>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARADDR>.
    //
    function automatic logic [((AXI_ADDRESS_WIDTH) - 1):0]   get_ARADDR(  );
        return ARADDR;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARADDR_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARADDR>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARADDR>.
    //
    function automatic logic   get_ARADDR_index1( int _this_dot_1 );
        return ARADDR[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARLEN
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARLEN>.
    //
    // Parameters:
    //     ARLEN_param - The value to set onto wire <ARLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLEN( logic [3:0] ARLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLEN = ARLEN_param;
        else
            m_ARLEN <= ARLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARLEN_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARLEN_param - The value to set onto wire <ARLEN>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLEN_index1( int _this_dot_1, logic  ARLEN_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLEN[_this_dot_1] = ARLEN_param;
        else
            m_ARLEN[_this_dot_1] <= ARLEN_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARLEN
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARLEN>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARLEN>.
    //
    function automatic logic [3:0]  get_ARLEN(  );
        return ARLEN;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARLEN_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARLEN>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARLEN>.
    //
    function automatic logic   get_ARLEN_index1( int _this_dot_1 );
        return ARLEN[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARSIZE
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARSIZE>.
    //
    // Parameters:
    //     ARSIZE_param - The value to set onto wire <ARSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARSIZE( logic [2:0] ARSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARSIZE = ARSIZE_param;
        else
            m_ARSIZE <= ARSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARSIZE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARSIZE_param - The value to set onto wire <ARSIZE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARSIZE_index1( int _this_dot_1, logic  ARSIZE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARSIZE[_this_dot_1] = ARSIZE_param;
        else
            m_ARSIZE[_this_dot_1] <= ARSIZE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARSIZE
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARSIZE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARSIZE>.
    //
    function automatic logic [2:0]  get_ARSIZE(  );
        return ARSIZE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARSIZE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARSIZE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARSIZE>.
    //
    function automatic logic   get_ARSIZE_index1( int _this_dot_1 );
        return ARSIZE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARBURST
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARBURST>.
    //
    // Parameters:
    //     ARBURST_param - The value to set onto wire <ARBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARBURST( logic [1:0] ARBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARBURST = ARBURST_param;
        else
            m_ARBURST <= ARBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARBURST_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARBURST_param - The value to set onto wire <ARBURST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARBURST_index1( int _this_dot_1, logic  ARBURST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARBURST[_this_dot_1] = ARBURST_param;
        else
            m_ARBURST[_this_dot_1] <= ARBURST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARBURST
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARBURST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARBURST>.
    //
    function automatic logic [1:0]  get_ARBURST(  );
        return ARBURST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARBURST_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARBURST>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARBURST>.
    //
    function automatic logic   get_ARBURST_index1( int _this_dot_1 );
        return ARBURST[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARLOCK
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARLOCK>.
    //
    // Parameters:
    //     ARLOCK_param - The value to set onto wire <ARLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLOCK( logic [1:0] ARLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLOCK = ARLOCK_param;
        else
            m_ARLOCK <= ARLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARLOCK_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARLOCK_param - The value to set onto wire <ARLOCK>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARLOCK_index1( int _this_dot_1, logic  ARLOCK_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARLOCK[_this_dot_1] = ARLOCK_param;
        else
            m_ARLOCK[_this_dot_1] <= ARLOCK_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARLOCK
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARLOCK>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARLOCK>.
    //
    function automatic logic [1:0]  get_ARLOCK(  );
        return ARLOCK;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARLOCK_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARLOCK>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARLOCK>.
    //
    function automatic logic   get_ARLOCK_index1( int _this_dot_1 );
        return ARLOCK[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARCACHE
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARCACHE>.
    //
    // Parameters:
    //     ARCACHE_param - The value to set onto wire <ARCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARCACHE( logic [3:0] ARCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARCACHE = ARCACHE_param;
        else
            m_ARCACHE <= ARCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARCACHE_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARCACHE_param - The value to set onto wire <ARCACHE>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARCACHE_index1( int _this_dot_1, logic  ARCACHE_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARCACHE[_this_dot_1] = ARCACHE_param;
        else
            m_ARCACHE[_this_dot_1] <= ARCACHE_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARCACHE
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARCACHE>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARCACHE>.
    //
    function automatic logic [3:0]  get_ARCACHE(  );
        return ARCACHE;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARCACHE_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARCACHE>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARCACHE>.
    //
    function automatic logic   get_ARCACHE_index1( int _this_dot_1 );
        return ARCACHE[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARPROT
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARPROT>.
    //
    // Parameters:
    //     ARPROT_param - The value to set onto wire <ARPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARPROT( logic [2:0] ARPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARPROT = ARPROT_param;
        else
            m_ARPROT <= ARPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARPROT_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARPROT_param - The value to set onto wire <ARPROT>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARPROT_index1( int _this_dot_1, logic  ARPROT_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARPROT[_this_dot_1] = ARPROT_param;
        else
            m_ARPROT[_this_dot_1] <= ARPROT_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARPROT
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARPROT>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARPROT>.
    //
    function automatic logic [2:0]  get_ARPROT(  );
        return ARPROT;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARPROT_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARPROT>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARPROT>.
    //
    function automatic logic   get_ARPROT_index1( int _this_dot_1 );
        return ARPROT[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARID
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARID>.
    //
    // Parameters:
    //     ARID_param - The value to set onto wire <ARID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARID( logic [((AXI_ID_WIDTH) - 1):0]  ARID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARID = ARID_param;
        else
            m_ARID <= ARID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARID_param - The value to set onto wire <ARID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARID_index1( int _this_dot_1, logic  ARID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARID[_this_dot_1] = ARID_param;
        else
            m_ARID[_this_dot_1] <= ARID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARID
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_ARID(  );
        return ARID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARID>.
    //
    function automatic logic   get_ARID_index1( int _this_dot_1 );
        return ARID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARREADY>.
    //
    // Parameters:
    //     ARREADY_param - The value to set onto wire <ARREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARREADY( logic ARREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARREADY = ARREADY_param;
        else
            m_ARREADY <= ARREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARREADY>.
    //
    function automatic logic get_ARREADY(  );
        return ARREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_ARUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <ARUSER>.
    //
    // Parameters:
    //     ARUSER_param - The value to set onto wire <ARUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARUSER( logic [7:0] ARUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARUSER = ARUSER_param;
        else
            m_ARUSER <= ARUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_ARUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <ARUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     ARUSER_param - The value to set onto wire <ARUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_ARUSER_index1( int _this_dot_1, logic  ARUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_ARUSER[_this_dot_1] = ARUSER_param;
        else
            m_ARUSER[_this_dot_1] <= ARUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_ARUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <ARUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <ARUSER>.
    //
    function automatic logic [7:0]  get_ARUSER(  );
        return ARUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_ARUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <ARUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <ARUSER>.
    //
    function automatic logic   get_ARUSER_index1( int _this_dot_1 );
        return ARUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <RVALID>.
    //
    // Parameters:
    //     RVALID_param - The value to set onto wire <RVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RVALID( logic RVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RVALID = RVALID_param;
        else
            m_RVALID <= RVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <RVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RVALID>.
    //
    function automatic logic get_RVALID(  );
        return RVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RLAST
    //-------------------------------------------------------------------------
    //     Set the value of wire <RLAST>.
    //
    // Parameters:
    //     RLAST_param - The value to set onto wire <RLAST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RLAST( logic RLAST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RLAST = RLAST_param;
        else
            m_RLAST <= RLAST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RLAST
    //-------------------------------------------------------------------------
    //     Get the value of wire <RLAST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RLAST>.
    //
    function automatic logic get_RLAST(  );
        return RLAST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RDATA
    //-------------------------------------------------------------------------
    //     Set the value of wire <RDATA>.
    //
    // Parameters:
    //     RDATA_param - The value to set onto wire <RDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RDATA( logic [((AXI_RDATA_WIDTH) - 1):0]  RDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RDATA = RDATA_param;
        else
            m_RDATA <= RDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RDATA_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RDATA_param - The value to set onto wire <RDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RDATA_index1( int _this_dot_1, logic  RDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RDATA[_this_dot_1] = RDATA_param;
        else
            m_RDATA[_this_dot_1] <= RDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RDATA
    //-------------------------------------------------------------------------
    //     Get the value of wire <RDATA>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RDATA>.
    //
    function automatic logic [((AXI_RDATA_WIDTH) - 1):0]   get_RDATA(  );
        return RDATA;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RDATA_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RDATA>.
    //
    function automatic logic   get_RDATA_index1( int _this_dot_1 );
        return RDATA[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RRESP
    //-------------------------------------------------------------------------
    //     Set the value of wire <RRESP>.
    //
    // Parameters:
    //     RRESP_param - The value to set onto wire <RRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RRESP( logic [1:0] RRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RRESP = RRESP_param;
        else
            m_RRESP <= RRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RRESP_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RRESP_param - The value to set onto wire <RRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RRESP_index1( int _this_dot_1, logic  RRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RRESP[_this_dot_1] = RRESP_param;
        else
            m_RRESP[_this_dot_1] <= RRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RRESP
    //-------------------------------------------------------------------------
    //     Get the value of wire <RRESP>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RRESP>.
    //
    function automatic logic [1:0]  get_RRESP(  );
        return RRESP;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RRESP_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RRESP>.
    //
    function automatic logic   get_RRESP_index1( int _this_dot_1 );
        return RRESP[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RID
    //-------------------------------------------------------------------------
    //     Set the value of wire <RID>.
    //
    // Parameters:
    //     RID_param - The value to set onto wire <RID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RID( logic [((AXI_ID_WIDTH) - 1):0]  RID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RID = RID_param;
        else
            m_RID <= RID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RID_param - The value to set onto wire <RID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RID_index1( int _this_dot_1, logic  RID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RID[_this_dot_1] = RID_param;
        else
            m_RID[_this_dot_1] <= RID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RID
    //-------------------------------------------------------------------------
    //     Get the value of wire <RID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_RID(  );
        return RID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RID>.
    //
    function automatic logic   get_RID_index1( int _this_dot_1 );
        return RID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <RREADY>.
    //
    // Parameters:
    //     RREADY_param - The value to set onto wire <RREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RREADY( logic RREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RREADY = RREADY_param;
        else
            m_RREADY <= RREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <RREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RREADY>.
    //
    function automatic logic get_RREADY(  );
        return RREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_RUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <RUSER>.
    //
    // Parameters:
    //     RUSER_param - The value to set onto wire <RUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RUSER( logic [7:0] RUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RUSER = RUSER_param;
        else
            m_RUSER <= RUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_RUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <RUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     RUSER_param - The value to set onto wire <RUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_RUSER_index1( int _this_dot_1, logic  RUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_RUSER[_this_dot_1] = RUSER_param;
        else
            m_RUSER[_this_dot_1] <= RUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_RUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <RUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <RUSER>.
    //
    function automatic logic [7:0]  get_RUSER(  );
        return RUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_RUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <RUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <RUSER>.
    //
    function automatic logic   get_RUSER_index1( int _this_dot_1 );
        return RUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <WVALID>.
    //
    // Parameters:
    //     WVALID_param - The value to set onto wire <WVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WVALID( logic WVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WVALID = WVALID_param;
        else
            m_WVALID <= WVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <WVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WVALID>.
    //
    function automatic logic get_WVALID(  );
        return WVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WLAST
    //-------------------------------------------------------------------------
    //     Set the value of wire <WLAST>.
    //
    // Parameters:
    //     WLAST_param - The value to set onto wire <WLAST>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WLAST( logic WLAST_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WLAST = WLAST_param;
        else
            m_WLAST <= WLAST_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WLAST
    //-------------------------------------------------------------------------
    //     Get the value of wire <WLAST>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WLAST>.
    //
    function automatic logic get_WLAST(  );
        return WLAST;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WDATA
    //-------------------------------------------------------------------------
    //     Set the value of wire <WDATA>.
    //
    // Parameters:
    //     WDATA_param - The value to set onto wire <WDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WDATA( logic [((AXI_WDATA_WIDTH) - 1):0]  WDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WDATA = WDATA_param;
        else
            m_WDATA <= WDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WDATA_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WDATA_param - The value to set onto wire <WDATA>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WDATA_index1( int _this_dot_1, logic  WDATA_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WDATA[_this_dot_1] = WDATA_param;
        else
            m_WDATA[_this_dot_1] <= WDATA_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WDATA
    //-------------------------------------------------------------------------
    //     Get the value of wire <WDATA>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WDATA>.
    //
    function automatic logic [((AXI_WDATA_WIDTH) - 1):0]   get_WDATA(  );
        return WDATA;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WDATA_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WDATA>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WDATA>.
    //
    function automatic logic   get_WDATA_index1( int _this_dot_1 );
        return WDATA[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WSTRB
    //-------------------------------------------------------------------------
    //     Set the value of wire <WSTRB>.
    //
    // Parameters:
    //     WSTRB_param - The value to set onto wire <WSTRB>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WSTRB( logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  WSTRB_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WSTRB = WSTRB_param;
        else
            m_WSTRB <= WSTRB_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WSTRB_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WSTRB>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WSTRB_param - The value to set onto wire <WSTRB>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WSTRB_index1( int _this_dot_1, logic  WSTRB_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WSTRB[_this_dot_1] = WSTRB_param;
        else
            m_WSTRB[_this_dot_1] <= WSTRB_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WSTRB
    //-------------------------------------------------------------------------
    //     Get the value of wire <WSTRB>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WSTRB>.
    //
    function automatic logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]   get_WSTRB(  );
        return WSTRB;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WSTRB_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WSTRB>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WSTRB>.
    //
    function automatic logic   get_WSTRB_index1( int _this_dot_1 );
        return WSTRB[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WID
    //-------------------------------------------------------------------------
    //     Set the value of wire <WID>.
    //
    // Parameters:
    //     WID_param - The value to set onto wire <WID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WID( logic [((AXI_ID_WIDTH) - 1):0]  WID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WID = WID_param;
        else
            m_WID <= WID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WID_param - The value to set onto wire <WID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WID_index1( int _this_dot_1, logic  WID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WID[_this_dot_1] = WID_param;
        else
            m_WID[_this_dot_1] <= WID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WID
    //-------------------------------------------------------------------------
    //     Get the value of wire <WID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_WID(  );
        return WID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WID>.
    //
    function automatic logic   get_WID_index1( int _this_dot_1 );
        return WID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <WREADY>.
    //
    // Parameters:
    //     WREADY_param - The value to set onto wire <WREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WREADY( logic WREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WREADY = WREADY_param;
        else
            m_WREADY <= WREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <WREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WREADY>.
    //
    function automatic logic get_WREADY(  );
        return WREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_WUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <WUSER>.
    //
    // Parameters:
    //     WUSER_param - The value to set onto wire <WUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WUSER( logic [7:0] WUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WUSER = WUSER_param;
        else
            m_WUSER <= WUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_WUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <WUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     WUSER_param - The value to set onto wire <WUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_WUSER_index1( int _this_dot_1, logic  WUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_WUSER[_this_dot_1] = WUSER_param;
        else
            m_WUSER[_this_dot_1] <= WUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_WUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <WUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <WUSER>.
    //
    function automatic logic [7:0]  get_WUSER(  );
        return WUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_WUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <WUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <WUSER>.
    //
    function automatic logic   get_WUSER_index1( int _this_dot_1 );
        return WUSER[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BVALID
    //-------------------------------------------------------------------------
    //     Set the value of wire <BVALID>.
    //
    // Parameters:
    //     BVALID_param - The value to set onto wire <BVALID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BVALID( logic BVALID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BVALID = BVALID_param;
        else
            m_BVALID <= BVALID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BVALID
    //-------------------------------------------------------------------------
    //     Get the value of wire <BVALID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BVALID>.
    //
    function automatic logic get_BVALID(  );
        return BVALID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BRESP
    //-------------------------------------------------------------------------
    //     Set the value of wire <BRESP>.
    //
    // Parameters:
    //     BRESP_param - The value to set onto wire <BRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BRESP( logic [1:0] BRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BRESP = BRESP_param;
        else
            m_BRESP <= BRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BRESP_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BRESP_param - The value to set onto wire <BRESP>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BRESP_index1( int _this_dot_1, logic  BRESP_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BRESP[_this_dot_1] = BRESP_param;
        else
            m_BRESP[_this_dot_1] <= BRESP_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BRESP
    //-------------------------------------------------------------------------
    //     Get the value of wire <BRESP>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BRESP>.
    //
    function automatic logic [1:0]  get_BRESP(  );
        return BRESP;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BRESP_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BRESP>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BRESP>.
    //
    function automatic logic   get_BRESP_index1( int _this_dot_1 );
        return BRESP[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BID
    //-------------------------------------------------------------------------
    //     Set the value of wire <BID>.
    //
    // Parameters:
    //     BID_param - The value to set onto wire <BID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BID( logic [((AXI_ID_WIDTH) - 1):0]  BID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BID = BID_param;
        else
            m_BID <= BID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BID_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BID_param - The value to set onto wire <BID>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BID_index1( int _this_dot_1, logic  BID_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BID[_this_dot_1] = BID_param;
        else
            m_BID[_this_dot_1] <= BID_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BID
    //-------------------------------------------------------------------------
    //     Get the value of wire <BID>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BID>.
    //
    function automatic logic [((AXI_ID_WIDTH) - 1):0]   get_BID(  );
        return BID;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BID_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BID>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BID>.
    //
    function automatic logic   get_BID_index1( int _this_dot_1 );
        return BID[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BREADY
    //-------------------------------------------------------------------------
    //     Set the value of wire <BREADY>.
    //
    // Parameters:
    //     BREADY_param - The value to set onto wire <BREADY>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BREADY( logic BREADY_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BREADY = BREADY_param;
        else
            m_BREADY <= BREADY_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BREADY
    //-------------------------------------------------------------------------
    //     Get the value of wire <BREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BREADY>.
    //
    function automatic logic get_BREADY(  );
        return BREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_BUSER
    //-------------------------------------------------------------------------
    //     Set the value of wire <BUSER>.
    //
    // Parameters:
    //     BUSER_param - The value to set onto wire <BUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BUSER( logic [7:0] BUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BUSER = BUSER_param;
        else
            m_BUSER <= BUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- set_BUSER_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of wire <BUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     BUSER_param - The value to set onto wire <BUSER>.
    //     non_blocking - Set to 1 for a non-blocking assignment.
    //
    task automatic set_BUSER_index1( int _this_dot_1, logic  BUSER_param = 'z, bit non_blocking = 1'b0 );
        if ( non_blocking == 1'b0 )
            m_BUSER[_this_dot_1] = BUSER_param;
        else
            m_BUSER[_this_dot_1] <= BUSER_param;
    endtask


    //-------------------------------------------------------------------------
    // Function:- get_BUSER
    //-------------------------------------------------------------------------
    //     Get the value of wire <BUSER>.
    //
    // Parameters:
    //
    // Returns the current value of the wire <BUSER>.
    //
    function automatic logic [7:0]  get_BUSER(  );
        return BUSER;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_BUSER_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of wire <BUSER>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the wire <BUSER>.
    //
    function automatic logic   get_BUSER_index1( int _this_dot_1 );
        return BUSER[_this_dot_1];
    endfunction

    //-------------------------------------------------------------------------
    // Tasks to wait for a change to a global variable with read access
    //-------------------------------------------------------------------------


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_write_ctrl_to_data_mintime
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_write_ctrl_to_data_mintime>.
    //
    task automatic wait_for_config_write_ctrl_to_data_mintime(  );
        begin
            @( config_write_ctrl_to_data_mintime );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_master_write_delay
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_master_write_delay>.
    //
    task automatic wait_for_config_master_write_delay(  );
        begin
            @( config_master_write_delay );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_all_assertions
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_all_assertions>.
    //
    task automatic wait_for_config_enable_all_assertions(  );
        begin
            @( config_enable_all_assertions );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_assertion
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_assertion>.
    //
    task automatic wait_for_config_enable_assertion(  );
        begin
            @( config_enable_assertion );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_enable_assertion_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_enable_assertion_index1( input int _this_dot_1 );
        begin
            @( config_enable_assertion[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_start_addr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_start_addr>.
    //
    task automatic wait_for_config_slave_start_addr(  );
        begin
            @( config_slave_start_addr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_start_addr_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_slave_start_addr_index1( input int _this_dot_1 );
        begin
            @( config_slave_start_addr[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_end_addr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_end_addr>.
    //
    task automatic wait_for_config_slave_end_addr(  );
        begin
            @( config_slave_end_addr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_slave_end_addr_index1
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    task automatic wait_for_config_slave_end_addr_index1( input int _this_dot_1 );
        begin
            @( config_slave_end_addr[_this_dot_1] );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_support_exclusive_access
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_support_exclusive_access>.
    //
    task automatic wait_for_config_support_exclusive_access(  );
        begin
            @( config_support_exclusive_access );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_read_data_reordering_depth
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_read_data_reordering_depth>.
    //
    task automatic wait_for_config_read_data_reordering_depth(  );
        begin
            @( config_read_data_reordering_depth );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_transaction_time_factor
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_transaction_time_factor>.
    //
    task automatic wait_for_config_max_transaction_time_factor(  );
        begin
            @( config_max_transaction_time_factor );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_timeout_max_data_transfer
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_timeout_max_data_transfer>.
    //
    task automatic wait_for_config_timeout_max_data_transfer(  );
        begin
            @( config_timeout_max_data_transfer );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_burst_timeout_factor
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_burst_timeout_factor>.
    //
    task automatic wait_for_config_burst_timeout_factor(  );
        begin
            @( config_burst_timeout_factor );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_AWVALID_assertion_to_AWREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    task automatic wait_for_config_max_latency_AWVALID_assertion_to_AWREADY(  );
        begin
            @( config_max_latency_AWVALID_assertion_to_AWREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_ARVALID_assertion_to_ARREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    task automatic wait_for_config_max_latency_ARVALID_assertion_to_ARREADY(  );
        begin
            @( config_max_latency_ARVALID_assertion_to_ARREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_RVALID_assertion_to_RREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_RVALID_assertion_to_RREADY>.
    //
    task automatic wait_for_config_max_latency_RVALID_assertion_to_RREADY(  );
        begin
            @( config_max_latency_RVALID_assertion_to_RREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_BVALID_assertion_to_BREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_BVALID_assertion_to_BREADY>.
    //
    task automatic wait_for_config_max_latency_BVALID_assertion_to_BREADY(  );
        begin
            @( config_max_latency_BVALID_assertion_to_BREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_latency_WVALID_assertion_to_WREADY
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_latency_WVALID_assertion_to_WREADY>.
    //
    task automatic wait_for_config_max_latency_WVALID_assertion_to_WREADY(  );
        begin
            @( config_max_latency_WVALID_assertion_to_WREADY );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_master_error_position
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_master_error_position>.
    //
    task automatic wait_for_config_master_error_position(  );
        begin
            @( config_master_error_position );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_setup_time
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_setup_time>.
    //
    task automatic wait_for_config_setup_time(  );
        begin
            @( config_setup_time );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_hold_time
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_hold_time>.
    //
    task automatic wait_for_config_hold_time(  );
        begin
            @( config_hold_time );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_wr
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_wr>.
    //
    task automatic wait_for_config_max_outstanding_wr(  );
        begin
            @( config_max_outstanding_wr );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_rd
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_rd>.
    //
    task automatic wait_for_config_max_outstanding_rd(  );
        begin
            @( config_max_outstanding_rd );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_max_outstanding_rw
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_max_outstanding_rw>.
    //
    task automatic wait_for_config_max_outstanding_rw(  );
        begin
            @( config_max_outstanding_rw );
        end
    endtask


    //------------------------------------------------------------------------------
    // Function:- wait_for_config_is_issuing
    //------------------------------------------------------------------------------
    //     Wait for a change on variable <axi::config_is_issuing>.
    //
    task automatic wait_for_config_is_issuing(  );
        begin
            @( config_is_issuing );
        end
    endtask


    //-------------------------------------------------------------------------
    // Functions to set global variables with write access
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- set_config_write_ctrl_to_data_mintime
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_write_ctrl_to_data_mintime>.
    //
    // Parameters:
    //     config_write_ctrl_to_data_mintime_param - The value to assign to variable <config_write_ctrl_to_data_mintime>.
    //
    function automatic void set_config_write_ctrl_to_data_mintime( int unsigned config_write_ctrl_to_data_mintime_param );
        config_write_ctrl_to_data_mintime = config_write_ctrl_to_data_mintime_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_master_write_delay
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_master_write_delay>.
    //
    // Parameters:
    //     config_master_write_delay_param - The value to assign to variable <config_master_write_delay>.
    //
    function automatic void set_config_master_write_delay( bit config_master_write_delay_param );
        config_master_write_delay = config_master_write_delay_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_all_assertions
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_enable_all_assertions>.
    //
    // Parameters:
    //     config_enable_all_assertions_param - The value to assign to variable <config_enable_all_assertions>.
    //
    function automatic void set_config_enable_all_assertions( bit config_enable_all_assertions_param );
        config_enable_all_assertions = config_enable_all_assertions_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_assertion
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_enable_assertion>.
    //
    // Parameters:
    //     config_enable_assertion_param - The value to assign to variable <config_enable_assertion>.
    //
    function automatic void set_config_enable_assertion( bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
        config_enable_assertion = config_enable_assertion_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_enable_assertion_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_enable_assertion_param - The value to assign to variable <config_enable_assertion>.
    //
    function automatic void set_config_enable_assertion_index1( int _this_dot_1, bit  config_enable_assertion_param );
        config_enable_assertion[_this_dot_1] = config_enable_assertion_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_start_addr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_slave_start_addr>.
    //
    // Parameters:
    //     config_slave_start_addr_param - The value to assign to variable <config_slave_start_addr>.
    //
    function automatic void set_config_slave_start_addr( bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param );
        config_slave_start_addr = config_slave_start_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_start_addr_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_slave_start_addr_param - The value to assign to variable <config_slave_start_addr>.
    //
    function automatic void set_config_slave_start_addr_index1( int _this_dot_1, bit  config_slave_start_addr_param );
        config_slave_start_addr[_this_dot_1] = config_slave_start_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_end_addr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_slave_end_addr>.
    //
    // Parameters:
    //     config_slave_end_addr_param - The value to assign to variable <config_slave_end_addr>.
    //
    function automatic void set_config_slave_end_addr( bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param );
        config_slave_end_addr = config_slave_end_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_slave_end_addr_index1
    //-------------------------------------------------------------------------
    //     Set the value of one element of variable <config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //     config_slave_end_addr_param - The value to assign to variable <config_slave_end_addr>.
    //
    function automatic void set_config_slave_end_addr_index1( int _this_dot_1, bit  config_slave_end_addr_param );
        config_slave_end_addr[_this_dot_1] = config_slave_end_addr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_support_exclusive_access
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_support_exclusive_access>.
    //
    // Parameters:
    //     config_support_exclusive_access_param - The value to assign to variable <config_support_exclusive_access>.
    //
    function automatic void set_config_support_exclusive_access( bit config_support_exclusive_access_param );
        config_support_exclusive_access = config_support_exclusive_access_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_read_data_reordering_depth
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_read_data_reordering_depth>.
    //
    // Parameters:
    //     config_read_data_reordering_depth_param - The value to assign to variable <config_read_data_reordering_depth>.
    //
    function automatic void set_config_read_data_reordering_depth( int unsigned config_read_data_reordering_depth_param );
        config_read_data_reordering_depth = config_read_data_reordering_depth_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_transaction_time_factor
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_transaction_time_factor>.
    //
    // Parameters:
    //     config_max_transaction_time_factor_param - The value to assign to variable <config_max_transaction_time_factor>.
    //
    function automatic void set_config_max_transaction_time_factor( int unsigned config_max_transaction_time_factor_param );
        config_max_transaction_time_factor = config_max_transaction_time_factor_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_timeout_max_data_transfer
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_timeout_max_data_transfer>.
    //
    // Parameters:
    //     config_timeout_max_data_transfer_param - The value to assign to variable <config_timeout_max_data_transfer>.
    //
    function automatic void set_config_timeout_max_data_transfer( int config_timeout_max_data_transfer_param );
        config_timeout_max_data_transfer = config_timeout_max_data_transfer_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_burst_timeout_factor
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_burst_timeout_factor>.
    //
    // Parameters:
    //     config_burst_timeout_factor_param - The value to assign to variable <config_burst_timeout_factor>.
    //
    function automatic void set_config_burst_timeout_factor( int unsigned config_burst_timeout_factor_param );
        config_burst_timeout_factor = config_burst_timeout_factor_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_AWVALID_assertion_to_AWREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    // Parameters:
    //     config_max_latency_AWVALID_assertion_to_AWREADY_param - The value to assign to variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    function automatic void set_config_max_latency_AWVALID_assertion_to_AWREADY( int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
        config_max_latency_AWVALID_assertion_to_AWREADY = config_max_latency_AWVALID_assertion_to_AWREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_ARVALID_assertion_to_ARREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    // Parameters:
    //     config_max_latency_ARVALID_assertion_to_ARREADY_param - The value to assign to variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    function automatic void set_config_max_latency_ARVALID_assertion_to_ARREADY( int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
        config_max_latency_ARVALID_assertion_to_ARREADY = config_max_latency_ARVALID_assertion_to_ARREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_RVALID_assertion_to_RREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    // Parameters:
    //     config_max_latency_RVALID_assertion_to_RREADY_param - The value to assign to variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    function automatic void set_config_max_latency_RVALID_assertion_to_RREADY( int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
        config_max_latency_RVALID_assertion_to_RREADY = config_max_latency_RVALID_assertion_to_RREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_BVALID_assertion_to_BREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    // Parameters:
    //     config_max_latency_BVALID_assertion_to_BREADY_param - The value to assign to variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    function automatic void set_config_max_latency_BVALID_assertion_to_BREADY( int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
        config_max_latency_BVALID_assertion_to_BREADY = config_max_latency_BVALID_assertion_to_BREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_latency_WVALID_assertion_to_WREADY
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    // Parameters:
    //     config_max_latency_WVALID_assertion_to_WREADY_param - The value to assign to variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    function automatic void set_config_max_latency_WVALID_assertion_to_WREADY( int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
        config_max_latency_WVALID_assertion_to_WREADY = config_max_latency_WVALID_assertion_to_WREADY_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_master_error_position
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_master_error_position>.
    //
    // Parameters:
    //     config_master_error_position_param - The value to assign to variable <config_master_error_position>.
    //
    function automatic void set_config_master_error_position( axi_error_e config_master_error_position_param );
        config_master_error_position = config_master_error_position_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_setup_time
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_setup_time>.
    //
    // Parameters:
    //     config_setup_time_param - The value to assign to variable <config_setup_time>.
    //
    function automatic void set_config_setup_time( int config_setup_time_param );
        config_setup_time = config_setup_time_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_hold_time
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_hold_time>.
    //
    // Parameters:
    //     config_hold_time_param - The value to assign to variable <config_hold_time>.
    //
    function automatic void set_config_hold_time( int config_hold_time_param );
        config_hold_time = config_hold_time_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_wr
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_wr>.
    //
    // Parameters:
    //     config_max_outstanding_wr_param - The value to assign to variable <config_max_outstanding_wr>.
    //
    function automatic void set_config_max_outstanding_wr( int config_max_outstanding_wr_param );
        config_max_outstanding_wr = config_max_outstanding_wr_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_rd
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_rd>.
    //
    // Parameters:
    //     config_max_outstanding_rd_param - The value to assign to variable <config_max_outstanding_rd>.
    //
    function automatic void set_config_max_outstanding_rd( int config_max_outstanding_rd_param );
        config_max_outstanding_rd = config_max_outstanding_rd_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_max_outstanding_rw
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_max_outstanding_rw>.
    //
    // Parameters:
    //     config_max_outstanding_rw_param - The value to assign to variable <config_max_outstanding_rw>.
    //
    function automatic void set_config_max_outstanding_rw( int config_max_outstanding_rw_param );
        config_max_outstanding_rw = config_max_outstanding_rw_param;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- set_config_is_issuing
    //-------------------------------------------------------------------------
    //     Set the value of variable <config_is_issuing>.
    //
    // Parameters:
    //     config_is_issuing_param - The value to assign to variable <config_is_issuing>.
    //
    function automatic void set_config_is_issuing( bit config_is_issuing_param );
        config_is_issuing = config_is_issuing_param;
    endfunction


    //-------------------------------------------------------------------------
    // Functions to get global variables with read access
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Function:- get_config_write_ctrl_to_data_mintime
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_write_ctrl_to_data_mintime>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_write_ctrl_to_data_mintime>.
    //
    function automatic int unsigned get_config_write_ctrl_to_data_mintime(  );
        return config_write_ctrl_to_data_mintime;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_master_write_delay
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_master_write_delay>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_master_write_delay>.
    //
    function automatic bit get_config_master_write_delay(  );
        axi_get_deprecated_config_master_write_delay_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_master_write_delay;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_all_assertions
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_enable_all_assertions>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_enable_all_assertions>.
    //
    function automatic bit get_config_enable_all_assertions(  );
        return config_enable_all_assertions;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_assertion
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_enable_assertion>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_enable_assertion>.
    //
    function automatic bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]   get_config_enable_assertion(  );
        return config_enable_assertion;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_enable_assertion_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_enable_assertion>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_enable_assertion>.
    //
    function automatic bit   get_config_enable_assertion_index1( int _this_dot_1 );
        return config_enable_assertion[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_start_addr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_slave_start_addr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_slave_start_addr>.
    //
    function automatic bit [((AXI_ADDRESS_WIDTH) - 1):0]   get_config_slave_start_addr(  );
        axi_get_deprecated_config_slave_start_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_start_addr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_start_addr_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_slave_start_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_slave_start_addr>.
    //
    function automatic bit   get_config_slave_start_addr_index1( int _this_dot_1 );
        axi_get_deprecated_config_slave_start_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_start_addr[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_end_addr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_slave_end_addr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_slave_end_addr>.
    //
    function automatic bit [((AXI_ADDRESS_WIDTH) - 1):0]   get_config_slave_end_addr(  );
        axi_get_deprecated_config_slave_end_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_end_addr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_slave_end_addr_index1
    //-------------------------------------------------------------------------
    //     Get the value of one element of variable <config_slave_end_addr>.
    //
    // Parameters:
    //    _this_dot_1 - The array index for dimension 1.
    //
    // Returns the current value of the variable <config_slave_end_addr>.
    //
    function automatic bit   get_config_slave_end_addr_index1( int _this_dot_1 );
        axi_get_deprecated_config_slave_end_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_slave_end_addr[_this_dot_1];
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_support_exclusive_access
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_support_exclusive_access>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_support_exclusive_access>.
    //
    function automatic bit get_config_support_exclusive_access(  );
        return config_support_exclusive_access;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_read_data_reordering_depth
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_read_data_reordering_depth>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_read_data_reordering_depth>.
    //
    function automatic int unsigned get_config_read_data_reordering_depth(  );
        return config_read_data_reordering_depth;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_transaction_time_factor
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_transaction_time_factor>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_transaction_time_factor>.
    //
    function automatic int unsigned get_config_max_transaction_time_factor(  );
        return config_max_transaction_time_factor;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_timeout_max_data_transfer
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_timeout_max_data_transfer>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_timeout_max_data_transfer>.
    //
    function automatic int get_config_timeout_max_data_transfer(  );
        return config_timeout_max_data_transfer;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_burst_timeout_factor
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_burst_timeout_factor>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_burst_timeout_factor>.
    //
    function automatic int unsigned get_config_burst_timeout_factor(  );
        return config_burst_timeout_factor;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_AWVALID_assertion_to_AWREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_AWVALID_assertion_to_AWREADY>.
    //
    function automatic int unsigned get_config_max_latency_AWVALID_assertion_to_AWREADY(  );
        return config_max_latency_AWVALID_assertion_to_AWREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_ARVALID_assertion_to_ARREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_ARVALID_assertion_to_ARREADY>.
    //
    function automatic int unsigned get_config_max_latency_ARVALID_assertion_to_ARREADY(  );
        return config_max_latency_ARVALID_assertion_to_ARREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_RVALID_assertion_to_RREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_RVALID_assertion_to_RREADY>.
    //
    function automatic int unsigned get_config_max_latency_RVALID_assertion_to_RREADY(  );
        return config_max_latency_RVALID_assertion_to_RREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_BVALID_assertion_to_BREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_BVALID_assertion_to_BREADY>.
    //
    function automatic int unsigned get_config_max_latency_BVALID_assertion_to_BREADY(  );
        return config_max_latency_BVALID_assertion_to_BREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_latency_WVALID_assertion_to_WREADY
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_latency_WVALID_assertion_to_WREADY>.
    //
    function automatic int unsigned get_config_max_latency_WVALID_assertion_to_WREADY(  );
        return config_max_latency_WVALID_assertion_to_WREADY;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_master_error_position
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_master_error_position>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_master_error_position>.
    //
    function automatic axi_error_e get_config_master_error_position(  );
        axi_get_deprecated_config_master_error_position_into_SystemVerilog( _interface_ref ); // DPI call to imported task
        return config_master_error_position;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_setup_time
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_setup_time>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_setup_time>.
    //
    function automatic int get_config_setup_time(  );
        return config_setup_time;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_hold_time
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_hold_time>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_hold_time>.
    //
    function automatic int get_config_hold_time(  );
        return config_hold_time;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_wr
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_wr>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_wr>.
    //
    function automatic int get_config_max_outstanding_wr(  );
        return config_max_outstanding_wr;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_rd
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_rd>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_rd>.
    //
    function automatic int get_config_max_outstanding_rd(  );
        return config_max_outstanding_rd;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_max_outstanding_rw
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_max_outstanding_rw>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_max_outstanding_rw>.
    //
    function automatic int get_config_max_outstanding_rw(  );
        return config_max_outstanding_rw;
    endfunction


    //-------------------------------------------------------------------------
    // Function:- get_config_is_issuing
    //-------------------------------------------------------------------------
    //     Get the value of variable <config_is_issuing>.
    //
    // Parameters:
    //
    // Returns the current value of the variable <config_is_issuing>.
    //
    function automatic bit get_config_is_issuing(  );
        return config_is_issuing;
    endfunction


    //-------------------------------------------------------------------------
    // Functions to set/get generic interface configuration
    //-------------------------------------------------------------------------

    function void set_interface
    (
        input int what = 0,
        input int arg1 = 0,
        input int arg2 = 0,
        input int arg3 = 0,
        input int arg4 = 0,
        input int arg5 = 0,
        input int arg6 = 0,
        input int arg7 = 0,
        input int arg8 = 0,
        input int arg9 = 0,
        input int arg10 = 0
    );
        axi_set_interface( what, arg1, arg2, arg3, arg4, arg5, arg6, arg7, arg8, arg9, arg10 );
    endfunction

    function int get_interface
    (
        input int what = 0,
        input int arg1 = 0,
        input int arg2 = 0,
        input int arg3 = 0,
        input int arg4 = 0,
        input int arg5 = 0,
        input int arg6 = 0,
        input int arg7 = 0,
        input int arg8 = 0,
        input int arg9 = 0
    );
        return axi_get_interface( what, arg1, arg2, arg3, arg4, arg5, arg6, arg7, arg8, arg9 );
    endfunction

    //-------------------------------------------------------------------------
    // Functions to get the hierarchic name of this interface
    //-------------------------------------------------------------------------
    function string get_full_name();
        return axi_get_full_name();
    endfunction

    //--------------------------------------------------------------------------
    //
    // Group:- Monitor Value Change on Variable
    //
    //--------------------------------------------------------------------------

    function automatic void axi_local_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( ref int unsigned config_write_ctrl_to_data_mintime_param );
            axi_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( _interface_ref,config_write_ctrl_to_data_mintime); // DPI call to imported task
        
            axi_propagate_config_write_ctrl_to_data_mintime_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_write_ctrl_to_data_mintime_from_SystemVerilog( config_write_ctrl_to_data_mintime );
            end
        end
    end

    function automatic void axi_local_set_config_master_write_delay_from_SystemVerilog( ref bit config_master_write_delay_param );
            axi_set_config_master_write_delay_from_SystemVerilog( _interface_ref,config_master_write_delay); // DPI call to imported task
        
            axi_propagate_config_master_write_delay_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_master_write_delay_from_SystemVerilog( config_master_write_delay );
            end
        end
    end

    function automatic void axi_local_set_config_enable_all_assertions_from_SystemVerilog( ref bit config_enable_all_assertions_param );
            axi_set_config_enable_all_assertions_from_SystemVerilog( _interface_ref,config_enable_all_assertions); // DPI call to imported task
        
            axi_propagate_config_enable_all_assertions_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_enable_all_assertions_from_SystemVerilog( config_enable_all_assertions );
            end
        end
    end

    function automatic void axi_local_set_config_enable_assertion_from_SystemVerilog( ref bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
            axi_set_config_enable_assertion_from_SystemVerilog( _interface_ref,config_enable_assertion); // DPI call to imported task
        
            axi_propagate_config_enable_assertion_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_enable_assertion_from_SystemVerilog( config_enable_assertion );
            end
        end
    end

    function automatic void axi_local_set_config_slave_start_addr_from_SystemVerilog( ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_start_addr_param );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ADDRESS_WIDTH ); _this_dot_1++)
        begin
            axi_set_config_slave_start_addr_from_SystemVerilog_index1( _interface_ref,_this_dot_1,config_slave_start_addr[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
            axi_propagate_config_slave_start_addr_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_slave_start_addr_from_SystemVerilog( config_slave_start_addr );
            end
        end
    end

    function automatic void axi_local_set_config_slave_end_addr_from_SystemVerilog( ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  config_slave_end_addr_param );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ADDRESS_WIDTH ); _this_dot_1++)
        begin
            axi_set_config_slave_end_addr_from_SystemVerilog_index1( _interface_ref,_this_dot_1,config_slave_end_addr[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
            axi_propagate_config_slave_end_addr_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_slave_end_addr_from_SystemVerilog( config_slave_end_addr );
            end
        end
    end

    function automatic void axi_local_set_config_support_exclusive_access_from_SystemVerilog( ref bit config_support_exclusive_access_param );
            axi_set_config_support_exclusive_access_from_SystemVerilog( _interface_ref,config_support_exclusive_access); // DPI call to imported task
        
            axi_propagate_config_support_exclusive_access_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_support_exclusive_access_from_SystemVerilog( config_support_exclusive_access );
            end
        end
    end

    function automatic void axi_local_set_config_read_data_reordering_depth_from_SystemVerilog( ref int unsigned config_read_data_reordering_depth_param );
            axi_set_config_read_data_reordering_depth_from_SystemVerilog( _interface_ref,config_read_data_reordering_depth); // DPI call to imported task
        
            axi_propagate_config_read_data_reordering_depth_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_read_data_reordering_depth_from_SystemVerilog( config_read_data_reordering_depth );
            end
        end
    end

    function automatic void axi_local_set_config_max_transaction_time_factor_from_SystemVerilog( ref int unsigned config_max_transaction_time_factor_param );
            axi_set_config_max_transaction_time_factor_from_SystemVerilog( _interface_ref,config_max_transaction_time_factor); // DPI call to imported task
        
            axi_propagate_config_max_transaction_time_factor_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_transaction_time_factor_from_SystemVerilog( config_max_transaction_time_factor );
            end
        end
    end

    function automatic void axi_local_set_config_timeout_max_data_transfer_from_SystemVerilog( ref int config_timeout_max_data_transfer_param );
            axi_set_config_timeout_max_data_transfer_from_SystemVerilog( _interface_ref,config_timeout_max_data_transfer); // DPI call to imported task
        
            axi_propagate_config_timeout_max_data_transfer_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_timeout_max_data_transfer_from_SystemVerilog( config_timeout_max_data_transfer );
            end
        end
    end

    function automatic void axi_local_set_config_burst_timeout_factor_from_SystemVerilog( ref int unsigned config_burst_timeout_factor_param );
            axi_set_config_burst_timeout_factor_from_SystemVerilog( _interface_ref,config_burst_timeout_factor); // DPI call to imported task
        
            axi_propagate_config_burst_timeout_factor_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_burst_timeout_factor_from_SystemVerilog( config_burst_timeout_factor );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( ref int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
            axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( _interface_ref,config_max_latency_AWVALID_assertion_to_AWREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog( config_max_latency_AWVALID_assertion_to_AWREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( ref int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
            axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( _interface_ref,config_max_latency_ARVALID_assertion_to_ARREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog( config_max_latency_ARVALID_assertion_to_ARREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( ref int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
            axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( _interface_ref,config_max_latency_RVALID_assertion_to_RREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog( config_max_latency_RVALID_assertion_to_RREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( ref int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
            axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( _interface_ref,config_max_latency_BVALID_assertion_to_BREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog( config_max_latency_BVALID_assertion_to_BREADY );
            end
        end
    end

    function automatic void axi_local_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( ref int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
            axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( _interface_ref,config_max_latency_WVALID_assertion_to_WREADY); // DPI call to imported task
        
            axi_propagate_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog( config_max_latency_WVALID_assertion_to_WREADY );
            end
        end
    end

    function automatic void axi_local_set_config_master_error_position_from_SystemVerilog( ref axi_error_e config_master_error_position_param );
            axi_set_config_master_error_position_from_SystemVerilog( _interface_ref,config_master_error_position); // DPI call to imported task
        
            axi_propagate_config_master_error_position_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_master_error_position_from_SystemVerilog( config_master_error_position );
            end
        end
    end

    function automatic void axi_local_set_config_setup_time_from_SystemVerilog( ref int config_setup_time_param );
            axi_set_config_setup_time_from_SystemVerilog( _interface_ref,config_setup_time); // DPI call to imported task
        
            axi_propagate_config_setup_time_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_setup_time_from_SystemVerilog( config_setup_time );
            end
        end
    end

    function automatic void axi_local_set_config_hold_time_from_SystemVerilog( ref int config_hold_time_param );
            axi_set_config_hold_time_from_SystemVerilog( _interface_ref,config_hold_time); // DPI call to imported task
        
            axi_propagate_config_hold_time_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_hold_time_from_SystemVerilog( config_hold_time );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_wr_from_SystemVerilog( ref int config_max_outstanding_wr_param );
            axi_set_config_max_outstanding_wr_from_SystemVerilog( _interface_ref,config_max_outstanding_wr); // DPI call to imported task
        
            axi_propagate_config_max_outstanding_wr_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_wr_from_SystemVerilog( config_max_outstanding_wr );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_rd_from_SystemVerilog( ref int config_max_outstanding_rd_param );
            axi_set_config_max_outstanding_rd_from_SystemVerilog( _interface_ref,config_max_outstanding_rd); // DPI call to imported task
        
            axi_propagate_config_max_outstanding_rd_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_rd_from_SystemVerilog( config_max_outstanding_rd );
            end
        end
    end

    function automatic void axi_local_set_config_max_outstanding_rw_from_SystemVerilog( ref int config_max_outstanding_rw_param );
            axi_set_config_max_outstanding_rw_from_SystemVerilog( _interface_ref,config_max_outstanding_rw); // DPI call to imported task
        
            axi_propagate_config_max_outstanding_rw_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_max_outstanding_rw_from_SystemVerilog( config_max_outstanding_rw );
            end
        end
    end

    function automatic void axi_local_set_config_is_issuing_from_SystemVerilog( ref bit config_is_issuing_param );
            axi_set_config_is_issuing_from_SystemVerilog( _interface_ref,config_is_issuing); // DPI call to imported task
        
            axi_propagate_config_is_issuing_from_SystemVerilog( _interface_ref ); // DPI call to imported task
    endfunction

    initial
    begin
        begin
            wait(_interface_ref != 0);
            forever
            begin
                @( * ) axi_local_set_config_is_issuing_from_SystemVerilog( config_is_issuing );
            end
        end
    end

    //-------------------------------------------------------------------------
    // Transaction interface
    //-------------------------------------------------------------------------

    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_rw_transaction_addr;
    function void axi_get_temp_static_rw_transaction_addr( input int _d1, output bit  _value );
        _value = temp_static_rw_transaction_addr[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_addr( input int _d1, input bit  _value );
        temp_static_rw_transaction_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_rw_transaction_id;
    function void axi_get_temp_static_rw_transaction_id( input int _d1, output bit  _value );
        _value = temp_static_rw_transaction_id[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_id( input int _d1, input bit  _value );
        temp_static_rw_transaction_id[_d1] = _value;
    endfunction
    bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] temp_static_rw_transaction_data_words [];
    function void axi_get_temp_static_rw_transaction_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_rw_transaction_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_rw_transaction_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_rw_transaction_data_words[_d1][_d2] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] temp_static_rw_transaction_write_strobes [];
    function void axi_get_temp_static_rw_transaction_write_strobes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_rw_transaction_write_strobes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_rw_transaction_write_strobes( input int _d1, input int _d2, input bit _value );
        temp_static_rw_transaction_write_strobes[_d1][_d2] = _value;
    endfunction
    axi_response_e temp_static_rw_transaction_resp[];
    function void axi_get_temp_static_rw_transaction_resp( input int _d1, output axi_response_e _value );
        _value = temp_static_rw_transaction_resp[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_resp( input int _d1, input axi_response_e _value );
        temp_static_rw_transaction_resp[_d1] = _value;
    endfunction
    bit [7:0] temp_static_rw_transaction_data_user [];
    function void axi_get_temp_static_rw_transaction_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_rw_transaction_data_user[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_rw_transaction_data_user[_d1] = _value;
    endfunction
    int temp_static_rw_transaction_write_data_beats_delay[];
    function void axi_get_temp_static_rw_transaction_write_data_beats_delay( input int _d1, output int _value );
        _value = temp_static_rw_transaction_write_data_beats_delay[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_write_data_beats_delay( input int _d1, input int _value );
        temp_static_rw_transaction_write_data_beats_delay[_d1] = _value;
    endfunction
    int temp_static_rw_transaction_data_valid_delay[];
    function void axi_get_temp_static_rw_transaction_data_valid_delay( input int _d1, output int _value );
        _value = temp_static_rw_transaction_data_valid_delay[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_data_valid_delay( input int _d1, input int _value );
        temp_static_rw_transaction_data_valid_delay[_d1] = _value;
    endfunction
    int temp_static_rw_transaction_data_ready_delay[];
    function void axi_get_temp_static_rw_transaction_data_ready_delay( input int _d1, output int _value );
        _value = temp_static_rw_transaction_data_ready_delay[_d1];
    endfunction
    function void axi_set_temp_static_rw_transaction_data_ready_delay( input int _d1, input int _value );
        temp_static_rw_transaction_data_ready_delay[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_AXI_read_addr;
    function void axi_get_temp_static_AXI_read_addr( input int _d1, output bit  _value );
        _value = temp_static_AXI_read_addr[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_addr( input int _d1, input bit  _value );
        temp_static_AXI_read_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_AXI_read_id;
    function void axi_get_temp_static_AXI_read_id( input int _d1, output bit  _value );
        _value = temp_static_AXI_read_id[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_id( input int _d1, input bit  _value );
        temp_static_AXI_read_id[_d1] = _value;
    endfunction
    bit [((AXI_RDATA_WIDTH) - 1):0] temp_static_AXI_read_data_words [];
    function void axi_get_temp_static_AXI_read_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_AXI_read_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_AXI_read_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_AXI_read_data_words[_d1][_d2] = _value;
    endfunction
    axi_response_e temp_static_AXI_read_resp[];
    function void axi_get_temp_static_AXI_read_resp( input int _d1, output axi_response_e _value );
        _value = temp_static_AXI_read_resp[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_resp( input int _d1, input axi_response_e _value );
        temp_static_AXI_read_resp[_d1] = _value;
    endfunction
    bit [7:0] temp_static_AXI_read_data_user [];
    function void axi_get_temp_static_AXI_read_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_AXI_read_data_user[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_AXI_read_data_user[_d1] = _value;
    endfunction
    longint temp_static_AXI_read_data_start_time[];
    function void axi_get_temp_static_AXI_read_data_start_time( input int _d1, output longint _value );
        _value = temp_static_AXI_read_data_start_time[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_data_start_time( input int _d1, input longint _value );
        temp_static_AXI_read_data_start_time[_d1] = _value;
    endfunction
    longint temp_static_AXI_read_data_end_time[];
    function void axi_get_temp_static_AXI_read_data_end_time( input int _d1, output longint _value );
        _value = temp_static_AXI_read_data_end_time[_d1];
    endfunction
    function void axi_set_temp_static_AXI_read_data_end_time( input int _d1, input longint _value );
        temp_static_AXI_read_data_end_time[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_AXI_write_addr;
    function void axi_get_temp_static_AXI_write_addr( input int _d1, output bit  _value );
        _value = temp_static_AXI_write_addr[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_addr( input int _d1, input bit  _value );
        temp_static_AXI_write_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_AXI_write_id;
    function void axi_get_temp_static_AXI_write_id( input int _d1, output bit  _value );
        _value = temp_static_AXI_write_id[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_id( input int _d1, input bit  _value );
        temp_static_AXI_write_id[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0] temp_static_AXI_write_data_words [];
    function void axi_get_temp_static_AXI_write_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_AXI_write_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_AXI_write_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_AXI_write_data_words[_d1][_d2] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] temp_static_AXI_write_write_strobes [];
    function void axi_get_temp_static_AXI_write_write_strobes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_AXI_write_write_strobes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_AXI_write_write_strobes( input int _d1, input int _d2, input bit _value );
        temp_static_AXI_write_write_strobes[_d1][_d2] = _value;
    endfunction
    bit [7:0] temp_static_AXI_write_data_user [];
    function void axi_get_temp_static_AXI_write_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_AXI_write_data_user[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_AXI_write_data_user[_d1] = _value;
    endfunction
    int temp_static_AXI_write_write_data_beats_delay[];
    function void axi_get_temp_static_AXI_write_write_data_beats_delay( input int _d1, output int _value );
        _value = temp_static_AXI_write_write_data_beats_delay[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_write_data_beats_delay( input int _d1, input int _value );
        temp_static_AXI_write_write_data_beats_delay[_d1] = _value;
    endfunction
    longint temp_static_AXI_write_data_start_time[];
    function void axi_get_temp_static_AXI_write_data_start_time( input int _d1, output longint _value );
        _value = temp_static_AXI_write_data_start_time[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_data_start_time( input int _d1, input longint _value );
        temp_static_AXI_write_data_start_time[_d1] = _value;
    endfunction
    longint temp_static_AXI_write_data_end_time[];
    function void axi_get_temp_static_AXI_write_data_end_time( input int _d1, output longint _value );
        _value = temp_static_AXI_write_data_end_time[_d1];
    endfunction
    function void axi_set_temp_static_AXI_write_data_end_time( input int _d1, input longint _value );
        temp_static_AXI_write_data_end_time[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0] temp_static_data_resp_data_words [];
    function void axi_get_temp_static_data_resp_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_data_resp_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_data_resp_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_data_resp_data_words[_d1][_d2] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] temp_static_data_resp_write_strobes [];
    function void axi_get_temp_static_data_resp_write_strobes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_data_resp_write_strobes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_data_resp_write_strobes( input int _d1, input int _d2, input bit _value );
        temp_static_data_resp_write_strobes[_d1][_d2] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_data_resp_id;
    function void axi_get_temp_static_data_resp_id( input int _d1, output bit  _value );
        _value = temp_static_data_resp_id[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_id( input int _d1, input bit  _value );
        temp_static_data_resp_id[_d1] = _value;
    endfunction
    bit [7:0] temp_static_data_resp_data_user [];
    function void axi_get_temp_static_data_resp_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_data_resp_data_user[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_data_resp_data_user[_d1] = _value;
    endfunction
    int temp_static_data_resp_write_data_beats_delay[];
    function void axi_get_temp_static_data_resp_write_data_beats_delay( input int _d1, output int _value );
        _value = temp_static_data_resp_write_data_beats_delay[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_write_data_beats_delay( input int _d1, input int _value );
        temp_static_data_resp_write_data_beats_delay[_d1] = _value;
    endfunction
    longint temp_static_data_resp_data_beat_start_time[];
    function void axi_get_temp_static_data_resp_data_beat_start_time( input int _d1, output longint _value );
        _value = temp_static_data_resp_data_beat_start_time[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_data_beat_start_time( input int _d1, input longint _value );
        temp_static_data_resp_data_beat_start_time[_d1] = _value;
    endfunction
    longint temp_static_data_resp_data_beat_end_time[];
    function void axi_get_temp_static_data_resp_data_beat_end_time( input int _d1, output longint _value );
        _value = temp_static_data_resp_data_beat_end_time[_d1];
    endfunction
    function void axi_set_temp_static_data_resp_data_beat_end_time( input int _d1, input longint _value );
        temp_static_data_resp_data_beat_end_time[_d1] = _value;
    endfunction
    bit [((AXI_RDATA_WIDTH) - 1):0] temp_static_read_data_burst_data_words [];
    function void axi_get_temp_static_read_data_burst_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_read_data_burst_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_read_data_burst_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_read_data_burst_data_words[_d1][_d2] = _value;
    endfunction
    axi_response_e temp_static_read_data_burst_resp[];
    function void axi_get_temp_static_read_data_burst_resp( input int _d1, output axi_response_e _value );
        _value = temp_static_read_data_burst_resp[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_resp( input int _d1, input axi_response_e _value );
        temp_static_read_data_burst_resp[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_data_burst_id;
    function void axi_get_temp_static_read_data_burst_id( input int _d1, output bit  _value );
        _value = temp_static_read_data_burst_id[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_id( input int _d1, input bit  _value );
        temp_static_read_data_burst_id[_d1] = _value;
    endfunction
    bit [7:0] temp_static_read_data_burst_data_user [];
    function void axi_get_temp_static_read_data_burst_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_read_data_burst_data_user[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_read_data_burst_data_user[_d1] = _value;
    endfunction
    longint temp_static_read_data_burst_data_start_time[];
    function void axi_get_temp_static_read_data_burst_data_start_time( input int _d1, output longint _value );
        _value = temp_static_read_data_burst_data_start_time[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_data_start_time( input int _d1, input longint _value );
        temp_static_read_data_burst_data_start_time[_d1] = _value;
    endfunction
    longint temp_static_read_data_burst_data_end_time[];
    function void axi_get_temp_static_read_data_burst_data_end_time( input int _d1, output longint _value );
        _value = temp_static_read_data_burst_data_end_time[_d1];
    endfunction
    function void axi_set_temp_static_read_data_burst_data_end_time( input int _d1, input longint _value );
        temp_static_read_data_burst_data_end_time[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0] temp_static_write_data_burst_data_words [];
    function void axi_get_temp_static_write_data_burst_data_words( input int _d1, input int _d2, output bit _value );
        _value = temp_static_write_data_burst_data_words[_d1][_d2];
    endfunction
    function void axi_set_temp_static_write_data_burst_data_words( input int _d1, input int _d2, input bit _value );
        temp_static_write_data_burst_data_words[_d1][_d2] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] temp_static_write_data_burst_write_strobes [];
    function void axi_get_temp_static_write_data_burst_write_strobes( input int _d1, input int _d2, output bit _value );
        _value = temp_static_write_data_burst_write_strobes[_d1][_d2];
    endfunction
    function void axi_set_temp_static_write_data_burst_write_strobes( input int _d1, input int _d2, input bit _value );
        temp_static_write_data_burst_write_strobes[_d1][_d2] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_data_burst_id;
    function void axi_get_temp_static_write_data_burst_id( input int _d1, output bit  _value );
        _value = temp_static_write_data_burst_id[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_id( input int _d1, input bit  _value );
        temp_static_write_data_burst_id[_d1] = _value;
    endfunction
    bit [7:0] temp_static_write_data_burst_data_user [];
    function void axi_get_temp_static_write_data_burst_data_user( input int _d1, output bit [7:0] _value  );
        _value = temp_static_write_data_burst_data_user[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_data_user( input int _d1, input bit [7:0] _value  );
        temp_static_write_data_burst_data_user[_d1] = _value;
    endfunction
    int temp_static_write_data_burst_write_data_beats_delay[];
    function void axi_get_temp_static_write_data_burst_write_data_beats_delay( input int _d1, output int _value );
        _value = temp_static_write_data_burst_write_data_beats_delay[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_write_data_beats_delay( input int _d1, input int _value );
        temp_static_write_data_burst_write_data_beats_delay[_d1] = _value;
    endfunction
    longint temp_static_write_data_burst_data_start_time[];
    function void axi_get_temp_static_write_data_burst_data_start_time( input int _d1, output longint _value );
        _value = temp_static_write_data_burst_data_start_time[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_data_start_time( input int _d1, input longint _value );
        temp_static_write_data_burst_data_start_time[_d1] = _value;
    endfunction
    longint temp_static_write_data_burst_data_end_time[];
    function void axi_get_temp_static_write_data_burst_data_end_time( input int _d1, output longint _value );
        _value = temp_static_write_data_burst_data_end_time[_d1];
    endfunction
    function void axi_set_temp_static_write_data_burst_data_end_time( input int _d1, input longint _value );
        temp_static_write_data_burst_data_end_time[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_read_addr_channel_phase_addr;
    function void axi_get_temp_static_read_addr_channel_phase_addr( input int _d1, output bit  _value );
        _value = temp_static_read_addr_channel_phase_addr[_d1];
    endfunction
    function void axi_set_temp_static_read_addr_channel_phase_addr( input int _d1, input bit  _value );
        temp_static_read_addr_channel_phase_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_addr_channel_phase_id;
    function void axi_get_temp_static_read_addr_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_read_addr_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_read_addr_channel_phase_id( input int _d1, input bit  _value );
        temp_static_read_addr_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_RDATA_WIDTH) - 1):0]  temp_static_read_channel_phase_data;
    function void axi_get_temp_static_read_channel_phase_data( input int _d1, output bit  _value );
        _value = temp_static_read_channel_phase_data[_d1];
    endfunction
    function void axi_set_temp_static_read_channel_phase_data( input int _d1, input bit  _value );
        temp_static_read_channel_phase_data[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_channel_phase_id;
    function void axi_get_temp_static_read_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_read_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_read_channel_phase_id( input int _d1, input bit  _value );
        temp_static_read_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_write_addr_channel_phase_addr;
    function void axi_get_temp_static_write_addr_channel_phase_addr( input int _d1, output bit  _value );
        _value = temp_static_write_addr_channel_phase_addr[_d1];
    endfunction
    function void axi_set_temp_static_write_addr_channel_phase_addr( input int _d1, input bit  _value );
        temp_static_write_addr_channel_phase_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_addr_channel_phase_id;
    function void axi_get_temp_static_write_addr_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_write_addr_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_write_addr_channel_phase_id( input int _d1, input bit  _value );
        temp_static_write_addr_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0]  temp_static_write_channel_phase_data;
    function void axi_get_temp_static_write_channel_phase_data( input int _d1, output bit  _value );
        _value = temp_static_write_channel_phase_data[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_phase_data( input int _d1, input bit  _value );
        temp_static_write_channel_phase_data[_d1] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  temp_static_write_channel_phase_write_strobes;
    function void axi_get_temp_static_write_channel_phase_write_strobes( input int _d1, output bit  _value );
        _value = temp_static_write_channel_phase_write_strobes[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_phase_write_strobes( input int _d1, input bit  _value );
        temp_static_write_channel_phase_write_strobes[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_channel_phase_id;
    function void axi_get_temp_static_write_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_write_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_phase_id( input int _d1, input bit  _value );
        temp_static_write_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_resp_channel_phase_id;
    function void axi_get_temp_static_write_resp_channel_phase_id( input int _d1, output bit  _value );
        _value = temp_static_write_resp_channel_phase_id[_d1];
    endfunction
    function void axi_set_temp_static_write_resp_channel_phase_id( input int _d1, input bit  _value );
        temp_static_write_resp_channel_phase_id[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_read_addr_channel_cycle_addr;
    function void axi_get_temp_static_read_addr_channel_cycle_addr( input int _d1, output bit  _value );
        _value = temp_static_read_addr_channel_cycle_addr[_d1];
    endfunction
    function void axi_set_temp_static_read_addr_channel_cycle_addr( input int _d1, input bit  _value );
        temp_static_read_addr_channel_cycle_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_addr_channel_cycle_id;
    function void axi_get_temp_static_read_addr_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_read_addr_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_read_addr_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_read_addr_channel_cycle_id[_d1] = _value;
    endfunction
    bit [((AXI_RDATA_WIDTH) - 1):0]  temp_static_read_channel_cycle_data;
    function void axi_get_temp_static_read_channel_cycle_data( input int _d1, output bit  _value );
        _value = temp_static_read_channel_cycle_data[_d1];
    endfunction
    function void axi_set_temp_static_read_channel_cycle_data( input int _d1, input bit  _value );
        temp_static_read_channel_cycle_data[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_read_channel_cycle_id;
    function void axi_get_temp_static_read_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_read_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_read_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_read_channel_cycle_id[_d1] = _value;
    endfunction
    bit [((AXI_ADDRESS_WIDTH) - 1):0]  temp_static_write_addr_channel_cycle_addr;
    function void axi_get_temp_static_write_addr_channel_cycle_addr( input int _d1, output bit  _value );
        _value = temp_static_write_addr_channel_cycle_addr[_d1];
    endfunction
    function void axi_set_temp_static_write_addr_channel_cycle_addr( input int _d1, input bit  _value );
        temp_static_write_addr_channel_cycle_addr[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_addr_channel_cycle_id;
    function void axi_get_temp_static_write_addr_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_write_addr_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_write_addr_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_write_addr_channel_cycle_id[_d1] = _value;
    endfunction
    bit [((AXI_WDATA_WIDTH) - 1):0]  temp_static_write_channel_cycle_data;
    function void axi_get_temp_static_write_channel_cycle_data( input int _d1, output bit  _value );
        _value = temp_static_write_channel_cycle_data[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_cycle_data( input int _d1, input bit  _value );
        temp_static_write_channel_cycle_data[_d1] = _value;
    endfunction
    bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  temp_static_write_channel_cycle_strb;
    function void axi_get_temp_static_write_channel_cycle_strb( input int _d1, output bit  _value );
        _value = temp_static_write_channel_cycle_strb[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_cycle_strb( input int _d1, input bit  _value );
        temp_static_write_channel_cycle_strb[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_channel_cycle_id;
    function void axi_get_temp_static_write_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_write_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_write_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_write_channel_cycle_id[_d1] = _value;
    endfunction
    bit [((AXI_ID_WIDTH) - 1):0]  temp_static_write_resp_channel_cycle_id;
    function void axi_get_temp_static_write_resp_channel_cycle_id( input int _d1, output bit  _value );
        _value = temp_static_write_resp_channel_cycle_id[_d1];
    endfunction
    function void axi_set_temp_static_write_resp_channel_cycle_id( input int _d1, input bit  _value );
        temp_static_write_resp_channel_cycle_id[_d1] = _value;
    endfunction
    task automatic dvc_activate_rw_transaction
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp[],
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref axi_rw_e read_or_write,
        ref int address_to_data_latency,
        ref int data_to_response_latency,
        ref int write_address_to_data_delay,
        ref int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        ref int address_valid_delay,
        ref int data_valid_delay[],
        ref int write_response_valid_delay,
        ref int address_ready_delay,
        ref int data_ready_delay[],
        ref int write_response_ready_delay,
        ref bit write_data_with_address,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_valid_delay_DIMS0;
                automatic int data_ready_delay_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_rw_transaction_addr = addr;
            temp_static_rw_transaction_id = id;
            data_words_DIMS0 = data_words.size();
            temp_static_rw_transaction_data_words = data_words;
            write_strobes_DIMS0 = write_strobes.size();
            temp_static_rw_transaction_write_strobes = write_strobes;
            resp_DIMS0 = resp.size();
            temp_static_rw_transaction_resp = resp;
            data_user_DIMS0 = data_user.size();
            temp_static_rw_transaction_data_user = data_user;
            write_data_beats_delay_DIMS0 = write_data_beats_delay.size();
            temp_static_rw_transaction_write_data_beats_delay = write_data_beats_delay;
            data_valid_delay_DIMS0 = data_valid_delay.size();
            temp_static_rw_transaction_data_valid_delay = data_valid_delay;
            data_ready_delay_DIMS0 = data_ready_delay.size();
            temp_static_rw_transaction_data_ready_delay = data_ready_delay;
            // Call function to provide sized params and ingoing unsized params sizes.
            // In addition gets back updated sizes of unsized params.
            axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, data_words_DIMS0, write_strobes_DIMS0, resp_DIMS0, addr_user, data_user_DIMS0, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay_DIMS0, address_valid_delay, data_valid_delay_DIMS0, write_response_valid_delay, address_ready_delay, data_ready_delay_DIMS0, write_response_ready_delay, write_data_with_address, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_rw_transaction_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_write_strobes.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_rw_transaction_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_write_data_beats_delay.delete();
            end
            if (data_valid_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_valid_delay = new [data_valid_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_valid_delay.delete();
            end
            if (data_ready_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_ready_delay = new [data_ready_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_ready_delay.delete();
            end
            // Call function to get the sized params
            axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, addr_user, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, address_valid_delay, write_response_valid_delay, address_ready_delay, write_response_ready_delay, write_data_with_address, _unit_id); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_rw_transaction_addr;
            id = temp_static_rw_transaction_id;
            data_words = temp_static_rw_transaction_data_words;
            temp_static_rw_transaction_data_words.delete();
            write_strobes = temp_static_rw_transaction_write_strobes;
            temp_static_rw_transaction_write_strobes.delete();
            resp = temp_static_rw_transaction_resp;
            temp_static_rw_transaction_resp.delete();
            data_user = temp_static_rw_transaction_data_user;
            temp_static_rw_transaction_data_user.delete();
            write_data_beats_delay = temp_static_rw_transaction_write_data_beats_delay;
            temp_static_rw_transaction_write_data_beats_delay.delete();
            data_valid_delay = temp_static_rw_transaction_data_valid_delay;
            temp_static_rw_transaction_data_valid_delay.delete();
            data_ready_delay = temp_static_rw_transaction_data_ready_delay;
            temp_static_rw_transaction_data_ready_delay.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_rw_transaction
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((((AXI_RDATA_WIDTH > AXI_WDATA_WIDTH) ? AXI_RDATA_WIDTH : AXI_WDATA_WIDTH)) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp[],
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output axi_rw_e read_or_write,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        output int address_valid_delay,
        ref int data_valid_delay[],
        output int write_response_valid_delay,
        output int address_ready_delay,
        ref int data_ready_delay[],
        output int write_response_ready_delay,
        output bit write_data_with_address,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_valid_delay_DIMS0;
                automatic int data_ready_delay_DIMS0;
            // Call function to get unsized params sizes.
            axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, resp_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_valid_delay_DIMS0, data_ready_delay_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_rw_transaction_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_write_strobes.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_rw_transaction_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_write_data_beats_delay.delete();
            end
            if (data_valid_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_valid_delay = new [data_valid_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_valid_delay.delete();
            end
            if (data_ready_delay_DIMS0 != 0)
            begin
                temp_static_rw_transaction_data_ready_delay = new [data_ready_delay_DIMS0];
            end
            else
            begin
                temp_static_rw_transaction_data_ready_delay.delete();
            end
            // Call function to get the sized params
            axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, addr_user, resp_user, read_or_write, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, address_valid_delay, write_response_valid_delay, address_ready_delay, write_response_ready_delay, write_data_with_address, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_rw_transaction_addr;
            id = temp_static_rw_transaction_id;
            data_words = temp_static_rw_transaction_data_words;
            temp_static_rw_transaction_data_words.delete();
            write_strobes = temp_static_rw_transaction_write_strobes;
            temp_static_rw_transaction_write_strobes.delete();
            resp = temp_static_rw_transaction_resp;
            temp_static_rw_transaction_resp.delete();
            data_user = temp_static_rw_transaction_data_user;
            temp_static_rw_transaction_data_user.delete();
            write_data_beats_delay = temp_static_rw_transaction_write_data_beats_delay;
            temp_static_rw_transaction_write_data_beats_delay.delete();
            data_valid_delay = temp_static_rw_transaction_data_valid_delay;
            temp_static_rw_transaction_data_valid_delay.delete();
            data_ready_delay = temp_static_rw_transaction_data_ready_delay;
            temp_static_rw_transaction_data_ready_delay.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_AXI_read
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref int address_to_data_latency,
        ref longint addr_start_time,
        ref longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        ref int address_valid_delay,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_AXI_read_addr = addr;
            temp_static_AXI_read_id = id;
            data_words_DIMS0 = data_words.size();
            temp_static_AXI_read_data_words = data_words;
            resp_DIMS0 = resp.size();
            temp_static_AXI_read_resp = resp;
            data_user_DIMS0 = data_user.size();
            temp_static_AXI_read_data_user = data_user;
            data_start_time_DIMS0 = data_start_time.size();
            temp_static_AXI_read_data_start_time = data_start_time;
            data_end_time_DIMS0 = data_end_time.size();
            temp_static_AXI_read_data_end_time = data_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            // In addition gets back updated sizes of unsized params.
            axi_AXI_read_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, data_words_DIMS0, resp_DIMS0, addr_user, data_user_DIMS0, address_to_data_latency, addr_start_time, addr_end_time, data_start_time_DIMS0, data_end_time_DIMS0, address_valid_delay, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_words.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_AXI_read_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_user.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, addr_user, address_to_data_latency, addr_start_time, addr_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_AXI_read_addr;
            id = temp_static_AXI_read_id;
            data_words = temp_static_AXI_read_data_words;
            temp_static_AXI_read_data_words.delete();
            resp = temp_static_AXI_read_resp;
            temp_static_AXI_read_resp.delete();
            data_user = temp_static_AXI_read_data_user;
            temp_static_AXI_read_data_user.delete();
            data_start_time = temp_static_AXI_read_data_start_time;
            temp_static_AXI_read_data_start_time.delete();
            data_end_time = temp_static_AXI_read_data_end_time;
            temp_static_AXI_read_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_AXI_read
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output int address_to_data_latency,
        output longint addr_start_time,
        output longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        output int address_valid_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_AXI_read_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, resp_DIMS0, data_user_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_words.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_AXI_read_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_user.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_AXI_read_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_read_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, addr_user, address_to_data_latency, addr_start_time, addr_end_time, address_valid_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_AXI_read_addr;
            id = temp_static_AXI_read_id;
            data_words = temp_static_AXI_read_data_words;
            temp_static_AXI_read_data_words.delete();
            resp = temp_static_AXI_read_resp;
            temp_static_AXI_read_resp.delete();
            data_user = temp_static_AXI_read_data_user;
            temp_static_AXI_read_data_user.delete();
            data_start_time = temp_static_AXI_read_data_start_time;
            temp_static_AXI_read_data_start_time.delete();
            data_end_time = temp_static_AXI_read_data_end_time;
            temp_static_AXI_read_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_AXI_write
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        ref axi_size_e size,
        ref axi_burst_e burst,
        ref axi_lock_e lock,
        ref axi_cache_e cache,
        ref axi_prot_e prot,
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [3:0] burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref axi_response_e resp,
        ref bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref int address_to_data_latency,
        ref int data_to_response_latency,
        ref int write_address_to_data_delay,
        ref int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        ref longint addr_start_time,
        ref longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        ref longint wr_resp_start_time,
        ref longint wr_resp_end_time,
        ref int address_valid_delay,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_AXI_write_addr = addr;
            temp_static_AXI_write_id = id;
            data_words_DIMS0 = data_words.size();
            temp_static_AXI_write_data_words = data_words;
            write_strobes_DIMS0 = write_strobes.size();
            temp_static_AXI_write_write_strobes = write_strobes;
            data_user_DIMS0 = data_user.size();
            temp_static_AXI_write_data_user = data_user;
            write_data_beats_delay_DIMS0 = write_data_beats_delay.size();
            temp_static_AXI_write_write_data_beats_delay = write_data_beats_delay;
            data_start_time_DIMS0 = data_start_time.size();
            temp_static_AXI_write_data_start_time = data_start_time;
            data_end_time_DIMS0 = data_end_time.size();
            temp_static_AXI_write_data_end_time = data_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            // In addition gets back updated sizes of unsized params.
            axi_AXI_write_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, data_words_DIMS0, write_strobes_DIMS0, resp, addr_user, data_user_DIMS0, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, write_data_beats_delay_DIMS0, addr_start_time, addr_end_time, data_start_time_DIMS0, data_end_time_DIMS0, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_AXI_write_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_AXI_write_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_write_data_beats_delay.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, resp, addr_user, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, addr_start_time, addr_end_time, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_AXI_write_addr;
            id = temp_static_AXI_write_id;
            data_words = temp_static_AXI_write_data_words;
            temp_static_AXI_write_data_words.delete();
            write_strobes = temp_static_AXI_write_write_strobes;
            temp_static_AXI_write_write_strobes.delete();
            data_user = temp_static_AXI_write_data_user;
            temp_static_AXI_write_data_user.delete();
            write_data_beats_delay = temp_static_AXI_write_write_data_beats_delay;
            temp_static_AXI_write_write_data_beats_delay.delete();
            data_start_time = temp_static_AXI_write_data_start_time;
            temp_static_AXI_write_data_start_time.delete();
            data_end_time = temp_static_AXI_write_data_end_time;
            temp_static_AXI_write_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_AXI_write
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [3:0] burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output axi_response_e resp,
        output bit [7:0] addr_user,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        ref int write_data_beats_delay[],
        output longint addr_start_time,
        output longint addr_end_time,
        ref longint data_start_time[],
        ref longint data_end_time[],
        output longint wr_resp_start_time,
        output longint wr_resp_end_time,
        output int address_valid_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_AXI_write_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_AXI_write_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_AXI_write_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_write_data_beats_delay.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_AXI_write_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_AXI_write_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, size, burst, lock, cache, prot, burst_length, resp, addr_user, resp_user, address_to_data_latency, data_to_response_latency, write_address_to_data_delay, write_data_to_address_delay, addr_start_time, addr_end_time, wr_resp_start_time, wr_resp_end_time, address_valid_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_AXI_write_addr;
            id = temp_static_AXI_write_id;
            data_words = temp_static_AXI_write_data_words;
            temp_static_AXI_write_data_words.delete();
            write_strobes = temp_static_AXI_write_write_strobes;
            temp_static_AXI_write_write_strobes.delete();
            data_user = temp_static_AXI_write_data_user;
            temp_static_AXI_write_data_user.delete();
            write_data_beats_delay = temp_static_AXI_write_write_data_beats_delay;
            temp_static_AXI_write_write_data_beats_delay.delete();
            data_start_time = temp_static_AXI_write_data_start_time;
            temp_static_AXI_write_data_start_time.delete();
            data_end_time = temp_static_AXI_write_data_end_time;
            temp_static_AXI_write_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_activate_data_resp
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        ref int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        ref bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref axi_response_e resp,
        ref bit [7:0] data_user [],
        ref bit [7:0] resp_user,
        ref longint data_start,
        ref longint data_end,
        ref longint response_start,
        ref int write_data_beats_delay[],
        ref longint data_beat_start_time[],
        ref longint data_beat_end_time[],
        ref longint response_end_time,
        input int _unit_id = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_beat_start_time_DIMS0;
                automatic int data_beat_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            data_words_DIMS0 = data_words.size();
            temp_static_data_resp_data_words = data_words;
            write_strobes_DIMS0 = write_strobes.size();
            temp_static_data_resp_write_strobes = write_strobes;
            temp_static_data_resp_id = id;
            data_user_DIMS0 = data_user.size();
            temp_static_data_resp_data_user = data_user;
            write_data_beats_delay_DIMS0 = write_data_beats_delay.size();
            temp_static_data_resp_write_data_beats_delay = write_data_beats_delay;
            data_beat_start_time_DIMS0 = data_beat_start_time.size();
            temp_static_data_resp_data_beat_start_time = data_beat_start_time;
            data_beat_end_time_DIMS0 = data_beat_end_time.size();
            temp_static_data_resp_data_beat_end_time = data_beat_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            // In addition gets back updated sizes of unsized params.
            axi_data_resp_ActivatesActivatingActivate_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, data_words_DIMS0, write_strobes_DIMS0, resp, data_user_DIMS0, resp_user, data_start, data_end, response_start, write_data_beats_delay_DIMS0, data_beat_start_time_DIMS0, data_beat_end_time_DIMS0, response_end_time, _unit_id); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_data_resp_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_data_resp_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_data_resp_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_data_resp_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_data_resp_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_data_resp_write_data_beats_delay.delete();
            end
            if (data_beat_start_time_DIMS0 != 0)
            begin
                temp_static_data_resp_data_beat_start_time = new [data_beat_start_time_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_beat_start_time.delete();
            end
            if (data_beat_end_time_DIMS0 != 0)
            begin
                temp_static_data_resp_data_beat_end_time = new [data_beat_end_time_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_beat_end_time.delete();
            end
            // Call function to get the sized params
            axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, resp, resp_user, data_start, data_end, response_start, response_end_time, _unit_id); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data_words = temp_static_data_resp_data_words;
            temp_static_data_resp_data_words.delete();
            write_strobes = temp_static_data_resp_write_strobes;
            temp_static_data_resp_write_strobes.delete();
            id = temp_static_data_resp_id;
            data_user = temp_static_data_resp_data_user;
            temp_static_data_resp_data_user.delete();
            write_data_beats_delay = temp_static_data_resp_write_data_beats_delay;
            temp_static_data_resp_write_data_beats_delay.delete();
            data_beat_start_time = temp_static_data_resp_data_beat_start_time;
            temp_static_data_resp_data_beat_start_time.delete();
            data_beat_end_time = temp_static_data_resp_data_beat_end_time;
            temp_static_data_resp_data_beat_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_data_resp
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output axi_response_e resp,
        ref bit [7:0] data_user [],
        output bit [7:0] resp_user,
        output longint data_start,
        output longint data_end,
        output longint response_start,
        ref int write_data_beats_delay[],
        ref longint data_beat_start_time[],
        ref longint data_beat_end_time[],
        output longint response_end_time,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_beat_start_time_DIMS0;
                automatic int data_beat_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_data_resp_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_beat_start_time_DIMS0, data_beat_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_data_resp_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_data_resp_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_data_resp_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_data_resp_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_data_resp_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_data_resp_write_data_beats_delay.delete();
            end
            if (data_beat_start_time_DIMS0 != 0)
            begin
                temp_static_data_resp_data_beat_start_time = new [data_beat_start_time_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_beat_start_time.delete();
            end
            if (data_beat_end_time_DIMS0 != 0)
            begin
                temp_static_data_resp_data_beat_end_time = new [data_beat_end_time_DIMS0];
            end
            else
            begin
                temp_static_data_resp_data_beat_end_time.delete();
            end
            // Call function to get the sized params
            axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, resp, resp_user, data_start, data_end, response_start, response_end_time, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data_words = temp_static_data_resp_data_words;
            temp_static_data_resp_data_words.delete();
            write_strobes = temp_static_data_resp_write_strobes;
            temp_static_data_resp_write_strobes.delete();
            id = temp_static_data_resp_id;
            data_user = temp_static_data_resp_data_user;
            temp_static_data_resp_data_user.delete();
            write_data_beats_delay = temp_static_data_resp_write_data_beats_delay;
            temp_static_data_resp_write_data_beats_delay.delete();
            data_beat_start_time = temp_static_data_resp_data_beat_start_time;
            temp_static_data_resp_data_beat_start_time.delete();
            data_beat_end_time = temp_static_data_resp_data_beat_end_time;
            temp_static_data_resp_data_beat_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            data_words_DIMS0 = data_words.size();
            temp_static_read_data_burst_data_words = data_words;
            resp_DIMS0 = resp.size();
            temp_static_read_data_burst_resp = resp;
            temp_static_read_data_burst_id = id;
            data_user_DIMS0 = data_user.size();
            temp_static_read_data_burst_data_user = data_user;
            data_start_time_DIMS0 = data_start_time.size();
            temp_static_read_data_burst_data_start_time = data_start_time;
            data_end_time_DIMS0 = data_end_time.size();
            temp_static_read_data_burst_data_end_time = data_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_data_burst_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, data_words_DIMS0, resp_DIMS0, data_user_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            temp_static_read_data_burst_data_words.delete();
            temp_static_read_data_burst_resp.delete();
            temp_static_read_data_burst_data_user.delete();
            temp_static_read_data_burst_data_start_time.delete();
            temp_static_read_data_burst_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [3:0] burst_length,
        ref bit [((AXI_RDATA_WIDTH) - 1):0] data_words [],
        ref axi_response_e resp[],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int resp_DIMS0;
                automatic int data_user_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, resp_DIMS0, data_user_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_read_data_burst_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_data_words.delete();
            end
            if (resp_DIMS0 != 0)
            begin
                temp_static_read_data_burst_resp = new [resp_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_resp.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_read_data_burst_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_data_user.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_read_data_burst_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_read_data_burst_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_read_data_burst_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data_words = temp_static_read_data_burst_data_words;
            temp_static_read_data_burst_data_words.delete();
            resp = temp_static_read_data_burst_resp;
            temp_static_read_data_burst_resp.delete();
            id = temp_static_read_data_burst_id;
            data_user = temp_static_read_data_burst_data_user;
            temp_static_read_data_burst_data_user.delete();
            data_start_time = temp_static_read_data_burst_data_start_time;
            temp_static_read_data_burst_data_start_time.delete();
            data_end_time = temp_static_read_data_burst_data_end_time;
            temp_static_read_data_burst_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref int write_data_beats_delay[],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            data_words_DIMS0 = data_words.size();
            temp_static_write_data_burst_data_words = data_words;
            write_strobes_DIMS0 = write_strobes.size();
            temp_static_write_data_burst_write_strobes = write_strobes;
            temp_static_write_data_burst_id = id;
            data_user_DIMS0 = data_user.size();
            temp_static_write_data_burst_data_user = data_user;
            write_data_beats_delay_DIMS0 = write_data_beats_delay.size();
            temp_static_write_data_burst_write_data_beats_delay = write_data_beats_delay;
            data_start_time_DIMS0 = data_start_time.size();
            temp_static_write_data_burst_data_start_time = data_start_time;
            data_end_time_DIMS0 = data_end_time.size();
            temp_static_write_data_burst_data_end_time = data_end_time;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_data_burst_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            temp_static_write_data_burst_data_words.delete();
            temp_static_write_data_burst_write_strobes.delete();
            temp_static_write_data_burst_data_user.delete();
            temp_static_write_data_burst_write_data_beats_delay.delete();
            temp_static_write_data_burst_data_start_time.delete();
            temp_static_write_data_burst_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_data_burst
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output int burst_length,
        ref bit [((AXI_WDATA_WIDTH) - 1):0] data_words [],
        ref bit [(((AXI_WDATA_WIDTH / 8)) - 1):0] write_strobes [],
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        ref bit [7:0] data_user [],
        ref int write_data_beats_delay[],
        ref longint data_start_time[],
        ref longint data_end_time[],
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
                automatic int data_words_DIMS0;
                automatic int write_strobes_DIMS0;
                automatic int data_user_DIMS0;
                automatic int write_data_beats_delay_DIMS0;
                automatic int data_start_time_DIMS0;
                automatic int data_end_time_DIMS0;
            // Call function to get unsized params sizes.
            axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, data_words_DIMS0, write_strobes_DIMS0, data_user_DIMS0, write_data_beats_delay_DIMS0, data_start_time_DIMS0, data_end_time_DIMS0, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            if (data_words_DIMS0 != 0)
            begin
                temp_static_write_data_burst_data_words = new [data_words_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_data_words.delete();
            end
            if (write_strobes_DIMS0 != 0)
            begin
                temp_static_write_data_burst_write_strobes = new [write_strobes_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_write_strobes.delete();
            end
            if (data_user_DIMS0 != 0)
            begin
                temp_static_write_data_burst_data_user = new [data_user_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_data_user.delete();
            end
            if (write_data_beats_delay_DIMS0 != 0)
            begin
                temp_static_write_data_burst_write_data_beats_delay = new [write_data_beats_delay_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_write_data_beats_delay.delete();
            end
            if (data_start_time_DIMS0 != 0)
            begin
                temp_static_write_data_burst_data_start_time = new [data_start_time_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_data_start_time.delete();
            end
            if (data_end_time_DIMS0 != 0)
            begin
                temp_static_write_data_burst_data_end_time = new [data_end_time_DIMS0];
            end
            else
            begin
                temp_static_write_data_burst_data_end_time.delete();
            end
            // Call function to get the sized params
            axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data_words = temp_static_write_data_burst_data_words;
            temp_static_write_data_burst_data_words.delete();
            write_strobes = temp_static_write_data_burst_write_strobes;
            temp_static_write_data_burst_write_strobes.delete();
            id = temp_static_write_data_burst_id;
            data_user = temp_static_write_data_burst_data_user;
            temp_static_write_data_burst_data_user.delete();
            write_data_beats_delay = temp_static_write_data_burst_write_data_beats_delay;
            temp_static_write_data_burst_write_data_beats_delay.delete();
            data_start_time = temp_static_write_data_burst_data_start_time;
            temp_static_write_data_burst_data_start_time.delete();
            data_end_time = temp_static_write_data_burst_data_end_time;
            temp_static_write_data_burst_data_end_time.delete();
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_read_addr_channel_phase_addr = addr;
            temp_static_read_addr_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_addr_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, size, burst, lock, cache, prot, addr_user, address_valid_delay, address_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_read_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, size, burst, lock, cache, prot, addr_user, address_valid_delay, address_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_read_addr_channel_phase_addr;
            id = temp_static_read_addr_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_read_channel_phase_data = data;
            temp_static_read_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, resp, data_user, data_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_read_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, last, resp, data_user, data_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data = temp_static_read_channel_phase_data;
            id = temp_static_read_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_addr_channel_phase_addr = addr;
            temp_static_write_addr_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_addr_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, size, burst, lock, cache, prot, addr_user, address_valid_delay, address_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_addr_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, size, burst, lock, cache, prot, addr_user, address_valid_delay, address_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_write_addr_channel_phase_addr;
            id = temp_static_write_addr_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_channel_phase_data = data;
            temp_static_write_channel_phase_write_strobes = write_strobes;
            temp_static_write_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, data_user, data_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  write_strobes,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        output int data_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, last, data_user, data_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data = temp_static_write_channel_phase_data;
            write_strobes = temp_static_write_channel_phase_write_strobes;
            id = temp_static_write_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_resp_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int write_response_ready_delay,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_resp_channel_phase_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_resp_channel_phase_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, resp, resp_user, write_response_ready_delay, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_resp_channel_phase
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        output int write_response_ready_delay,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_resp_channel_phase_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, resp, resp_user, write_response_ready_delay, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            id = temp_static_write_resp_channel_phase_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_read_addr_channel_cycle_addr = addr;
            temp_static_read_addr_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, size, burst, lock, cache, prot, addr_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_read_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, size, burst, lock, cache, prot, addr_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_read_addr_channel_cycle_addr;
            id = temp_static_read_addr_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_read_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_read_channel_cycle_data = data;
            temp_static_read_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_read_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, resp, data_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_read_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_RDATA_WIDTH) - 1):0]  data,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_read_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, last, resp, data_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data = temp_static_read_channel_cycle_data;
            id = temp_static_read_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_read_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_read_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] addr_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_addr_channel_cycle_addr = addr;
            temp_static_write_addr_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, burst_length, size, burst, lock, cache, prot, addr_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_addr_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit [((AXI_ADDRESS_WIDTH) - 1):0]  addr,
        output bit [3:0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] addr_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, burst_length, size, burst, lock, cache, prot, addr_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            addr = temp_static_write_addr_channel_cycle_addr;
            id = temp_static_write_addr_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_addr_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        input bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] data_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_channel_cycle_data = data;
            temp_static_write_channel_cycle_strb = strb;
            temp_static_write_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, last, data_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit last,
        output bit [((AXI_WDATA_WIDTH) - 1):0]  data,
        output bit [(((AXI_WDATA_WIDTH / 8)) - 1):0]  strb,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] data_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, last, data_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            data = temp_static_write_channel_cycle_data;
            strb = temp_static_write_channel_cycle_strb;
            id = temp_static_write_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask

    task automatic dvc_put_write_resp_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [((AXI_ID_WIDTH) - 1):0]  id,
        input bit [7:0] resp_user,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Pass to CY the size of each open dimension (assumes rectangular arrays)
            // In addition copy any unsized or flexibly sized parameters to a related static variable which will be accessed element by element from the C
            temp_static_write_resp_channel_cycle_id = id;
            // Call function to provide sized params and ingoing unsized params sizes.
            axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, resp, resp_user, _unit_id); // DPI call to imported task
            // Delete the storage allocated for the static variable(s)
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_get_write_resp_channel_cycle
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output axi_response_e resp,
        output bit [((AXI_ID_WIDTH) - 1):0]  id,
        output bit [7:0] resp_user,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin
            int _trans_id;

            wait(_interface_ref != 0);

            // the real code .....
            // Create an array to hold the unsized dims for each param (..._DIMS)
            begin // Block to create unsized data arrays
            // Call function to get unsized params sizes.
            axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, _trans_id, _unit_id, _using); // DPI call to imported task
            // Create each unsized param
            // Call function to get the sized params
            axi_write_resp_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog(_comms_semantic,_as_end, _trans_id, resp, resp_user, _unit_id, _using); // DPI call to imported task
            // Copy unsized data from static variable(s) which has/have been set element by element from the C++
            // In addition delete the storage allocated for the static variable(s)
            id = temp_static_write_resp_channel_cycle_id;
            end // Block to create unsized data arrays
        end
    endtask

    task automatic dvc_put_write_resp_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_ready_SendSendingSent_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id); // DPI call to imported task
        end
    endtask

    task automatic dvc_get_write_resp_channel_ready
    (
        input questa_mvc_item_comms_semantic _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id = 0,
        input bit _using = 0
    );
        begin

            wait(_interface_ref != 0);

            // the real code .....
            // Call function to set/get the params, all are of known size
            axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog(_comms_semantic,_as_end, ready, _unit_id, _using); // DPI call to imported task
        end
    endtask


    //-------------------------------------------------------------------------
    // Generic Interface Configuration Support
    //

    import "DPI-C" context axi_set_interface = function void axi_set_interface
    (
        input int what,
        input int arg1,
        input int arg2,
        input int arg3,
        input int arg4,
        input int arg5,
        input int arg6,
        input int arg7,
        input int arg8,
        input int arg9,
        input int arg10
    );
    import "DPI-C" context axi_get_interface = function int axi_get_interface
    (
        input int what,
        input int arg1,
        input int arg2,
        input int arg3,
        input int arg4,
        input int arg5,
        input int arg6,
        input int arg7,
        input int arg8,
        input int arg9
    );


    //-------------------------------------------------------------------------
    // Functions to get the hierarchic name of this interface
    //
    import "DPI-C" context axi_get_full_name = function string axi_get_full_name();


    //-------------------------------------------------------------------------
    // Abstraction level Support
    //

    import "DPI-C" context axi_set_master_end_abstraction_level =
    function void axi_set_master_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_master_end_abstraction_level =
    function void axi_get_master_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_slave_end_abstraction_level =
    function void axi_set_slave_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_slave_end_abstraction_level =
    function void axi_get_slave_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_clock_source_end_abstraction_level =
    function void axi_set_clock_source_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_clock_source_end_abstraction_level =
    function void axi_get_clock_source_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );
    import "DPI-C" context axi_set_reset_source_end_abstraction_level =
    function void axi_set_reset_source_end_abstraction_level
    (
        input bit         wire_level,
        input bit         TLM_level
    );
    import "DPI-C" context axi_get_reset_source_end_abstraction_level =
    function void axi_get_reset_source_end_abstraction_level
    (
        output bit         wire_level,
        output bit         TLM_level
    );

    //-------------------------------------------------------------------------
    // Wire Level Interface Support
    //
    logic internal_ACLK = 'z;
    logic internal_ARESETn = 'z;
    logic internal_AWVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  internal_AWADDR = 'z;
    logic [3:0] internal_AWLEN = 'z;
    logic [2:0] internal_AWSIZE = 'z;
    logic [1:0] internal_AWBURST = 'z;
    logic [1:0] internal_AWLOCK = 'z;
    logic [3:0] internal_AWCACHE = 'z;
    logic [2:0] internal_AWPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_AWID = 'z;
    logic internal_AWREADY = 'z;
    logic [7:0] internal_AWUSER = 'z;
    logic internal_ARVALID = 'z;
    logic [((AXI_ADDRESS_WIDTH) - 1):0]  internal_ARADDR = 'z;
    logic [3:0] internal_ARLEN = 'z;
    logic [2:0] internal_ARSIZE = 'z;
    logic [1:0] internal_ARBURST = 'z;
    logic [1:0] internal_ARLOCK = 'z;
    logic [3:0] internal_ARCACHE = 'z;
    logic [2:0] internal_ARPROT = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_ARID = 'z;
    logic internal_ARREADY = 'z;
    logic [7:0] internal_ARUSER = 'z;
    logic internal_RVALID = 'z;
    logic internal_RLAST = 'z;
    logic [((AXI_RDATA_WIDTH) - 1):0]  internal_RDATA = 'z;
    logic [1:0] internal_RRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_RID = 'z;
    logic internal_RREADY = 'z;
    logic [7:0] internal_RUSER = 'z;
    logic internal_WVALID = 'z;
    logic internal_WLAST = 'z;
    logic [((AXI_WDATA_WIDTH) - 1):0]  internal_WDATA = 'z;
    logic [(((AXI_WDATA_WIDTH / 8)) - 1):0]  internal_WSTRB = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_WID = 'z;
    logic internal_WREADY = 'z;
    logic [7:0] internal_WUSER = 'z;
    logic internal_BVALID = 'z;
    logic [1:0] internal_BRESP = 'z;
    logic [((AXI_ID_WIDTH) - 1):0]  internal_BID = 'z;
    logic internal_BREADY = 'z;
    logic [7:0] internal_BUSER = 'z;

    import "DPI-C" context function void axi_set_ACLK_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit ACLK_param
    );
    import "DPI-C" context function void axi_propagate_ACLK_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ACLK_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit ACLK_param

    );
    export "DPI-C" function axi_initialise_ACLK_from_CY;

    import "DPI-C" context function void axi_set_ARESETn_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARESETn_param
    );
    import "DPI-C" context function void axi_propagate_ARESETn_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARESETn_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARESETn_param

    );
    export "DPI-C" function axi_initialise_ARESETn_from_CY;

    import "DPI-C" context function void axi_set_AWVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic AWVALID_param
    );
    import "DPI-C" context function void axi_propagate_AWVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic AWVALID_param

    );
    export "DPI-C" function axi_initialise_AWVALID_from_CY;

    import "DPI-C" context function void axi_set_AWADDR_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  AWADDR_param
    );
    import "DPI-C" context function void axi_propagate_AWADDR_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWADDR_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_AWADDR_from_CY_index1;
    export "DPI-C" function axi_initialise_AWADDR_from_CY;

    import "DPI-C" context function void axi_set_AWLEN_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] AWLEN_param
    );
    import "DPI-C" context function void axi_propagate_AWLEN_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWLEN_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] AWLEN_param

    );
    export "DPI-C" function axi_initialise_AWLEN_from_CY;

    import "DPI-C" context function void axi_set_AWSIZE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] AWSIZE_param
    );
    import "DPI-C" context function void axi_propagate_AWSIZE_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWSIZE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] AWSIZE_param

    );
    export "DPI-C" function axi_initialise_AWSIZE_from_CY;

    import "DPI-C" context function void axi_set_AWBURST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] AWBURST_param
    );
    import "DPI-C" context function void axi_propagate_AWBURST_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWBURST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] AWBURST_param

    );
    export "DPI-C" function axi_initialise_AWBURST_from_CY;

    import "DPI-C" context function void axi_set_AWLOCK_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] AWLOCK_param
    );
    import "DPI-C" context function void axi_propagate_AWLOCK_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWLOCK_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] AWLOCK_param

    );
    export "DPI-C" function axi_initialise_AWLOCK_from_CY;

    import "DPI-C" context function void axi_set_AWCACHE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] AWCACHE_param
    );
    import "DPI-C" context function void axi_propagate_AWCACHE_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWCACHE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] AWCACHE_param

    );
    export "DPI-C" function axi_initialise_AWCACHE_from_CY;

    import "DPI-C" context function void axi_set_AWPROT_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] AWPROT_param
    );
    import "DPI-C" context function void axi_propagate_AWPROT_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWPROT_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] AWPROT_param

    );
    export "DPI-C" function axi_initialise_AWPROT_from_CY;

    import "DPI-C" context function void axi_set_AWID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  AWID_param
    );
    import "DPI-C" context function void axi_propagate_AWID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_AWID_from_CY_index1;
    export "DPI-C" function axi_initialise_AWID_from_CY;

    import "DPI-C" context function void axi_set_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic AWREADY_param
    );
    import "DPI-C" context function void axi_propagate_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic AWREADY_param

    );
    export "DPI-C" function axi_initialise_AWREADY_from_CY;

    import "DPI-C" context function void axi_set_AWUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] AWUSER_param
    );
    import "DPI-C" context function void axi_propagate_AWUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_AWUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] AWUSER_param

    );
    export "DPI-C" function axi_initialise_AWUSER_from_CY;

    import "DPI-C" context function void axi_set_ARVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARVALID_param
    );
    import "DPI-C" context function void axi_propagate_ARVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARVALID_param

    );
    export "DPI-C" function axi_initialise_ARVALID_from_CY;

    import "DPI-C" context function void axi_set_ARADDR_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  ARADDR_param
    );
    import "DPI-C" context function void axi_propagate_ARADDR_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARADDR_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_ARADDR_from_CY_index1;
    export "DPI-C" function axi_initialise_ARADDR_from_CY;

    import "DPI-C" context function void axi_set_ARLEN_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] ARLEN_param
    );
    import "DPI-C" context function void axi_propagate_ARLEN_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARLEN_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] ARLEN_param

    );
    export "DPI-C" function axi_initialise_ARLEN_from_CY;

    import "DPI-C" context function void axi_set_ARSIZE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] ARSIZE_param
    );
    import "DPI-C" context function void axi_propagate_ARSIZE_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARSIZE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] ARSIZE_param

    );
    export "DPI-C" function axi_initialise_ARSIZE_from_CY;

    import "DPI-C" context function void axi_set_ARBURST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] ARBURST_param
    );
    import "DPI-C" context function void axi_propagate_ARBURST_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARBURST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] ARBURST_param

    );
    export "DPI-C" function axi_initialise_ARBURST_from_CY;

    import "DPI-C" context function void axi_set_ARLOCK_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] ARLOCK_param
    );
    import "DPI-C" context function void axi_propagate_ARLOCK_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARLOCK_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] ARLOCK_param

    );
    export "DPI-C" function axi_initialise_ARLOCK_from_CY;

    import "DPI-C" context function void axi_set_ARCACHE_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [3:0] ARCACHE_param
    );
    import "DPI-C" context function void axi_propagate_ARCACHE_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARCACHE_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [3:0] ARCACHE_param

    );
    export "DPI-C" function axi_initialise_ARCACHE_from_CY;

    import "DPI-C" context function void axi_set_ARPROT_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [2:0] ARPROT_param
    );
    import "DPI-C" context function void axi_propagate_ARPROT_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARPROT_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [2:0] ARPROT_param

    );
    export "DPI-C" function axi_initialise_ARPROT_from_CY;

    import "DPI-C" context function void axi_set_ARID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  ARID_param
    );
    import "DPI-C" context function void axi_propagate_ARID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_ARID_from_CY_index1;
    export "DPI-C" function axi_initialise_ARID_from_CY;

    import "DPI-C" context function void axi_set_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic ARREADY_param
    );
    import "DPI-C" context function void axi_propagate_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic ARREADY_param

    );
    export "DPI-C" function axi_initialise_ARREADY_from_CY;

    import "DPI-C" context function void axi_set_ARUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] ARUSER_param
    );
    import "DPI-C" context function void axi_propagate_ARUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_ARUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] ARUSER_param

    );
    export "DPI-C" function axi_initialise_ARUSER_from_CY;

    import "DPI-C" context function void axi_set_RVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RVALID_param
    );
    import "DPI-C" context function void axi_propagate_RVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RVALID_param

    );
    export "DPI-C" function axi_initialise_RVALID_from_CY;

    import "DPI-C" context function void axi_set_RLAST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RLAST_param
    );
    import "DPI-C" context function void axi_propagate_RLAST_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RLAST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RLAST_param

    );
    export "DPI-C" function axi_initialise_RLAST_from_CY;

    import "DPI-C" context function void axi_set_RDATA_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  RDATA_param
    );
    import "DPI-C" context function void axi_propagate_RDATA_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RDATA_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_RDATA_from_CY_index1;
    export "DPI-C" function axi_initialise_RDATA_from_CY;

    import "DPI-C" context function void axi_set_RRESP_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] RRESP_param
    );
    import "DPI-C" context function void axi_propagate_RRESP_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RRESP_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] RRESP_param

    );
    export "DPI-C" function axi_initialise_RRESP_from_CY;

    import "DPI-C" context function void axi_set_RID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  RID_param
    );
    import "DPI-C" context function void axi_propagate_RID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_RID_from_CY_index1;
    export "DPI-C" function axi_initialise_RID_from_CY;

    import "DPI-C" context function void axi_set_RREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic RREADY_param
    );
    import "DPI-C" context function void axi_propagate_RREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic RREADY_param

    );
    export "DPI-C" function axi_initialise_RREADY_from_CY;

    import "DPI-C" context function void axi_set_RUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] RUSER_param
    );
    import "DPI-C" context function void axi_propagate_RUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_RUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] RUSER_param

    );
    export "DPI-C" function axi_initialise_RUSER_from_CY;

    import "DPI-C" context function void axi_set_WVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WVALID_param
    );
    import "DPI-C" context function void axi_propagate_WVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WVALID_param

    );
    export "DPI-C" function axi_initialise_WVALID_from_CY;

    import "DPI-C" context function void axi_set_WLAST_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WLAST_param
    );
    import "DPI-C" context function void axi_propagate_WLAST_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WLAST_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WLAST_param

    );
    export "DPI-C" function axi_initialise_WLAST_from_CY;

    import "DPI-C" context function void axi_set_WDATA_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  WDATA_param
    );
    import "DPI-C" context function void axi_propagate_WDATA_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WDATA_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_WDATA_from_CY_index1;
    export "DPI-C" function axi_initialise_WDATA_from_CY;

    import "DPI-C" context function void axi_set_WSTRB_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  WSTRB_param
    );
    import "DPI-C" context function void axi_propagate_WSTRB_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WSTRB_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_WSTRB_from_CY_index1;
    export "DPI-C" function axi_initialise_WSTRB_from_CY;

    import "DPI-C" context function void axi_set_WID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  WID_param
    );
    import "DPI-C" context function void axi_propagate_WID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_WID_from_CY_index1;
    export "DPI-C" function axi_initialise_WID_from_CY;

    import "DPI-C" context function void axi_set_WREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic WREADY_param
    );
    import "DPI-C" context function void axi_propagate_WREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic WREADY_param

    );
    export "DPI-C" function axi_initialise_WREADY_from_CY;

    import "DPI-C" context function void axi_set_WUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] WUSER_param
    );
    import "DPI-C" context function void axi_propagate_WUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_WUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] WUSER_param

    );
    export "DPI-C" function axi_initialise_WUSER_from_CY;

    import "DPI-C" context function void axi_set_BVALID_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic BVALID_param
    );
    import "DPI-C" context function void axi_propagate_BVALID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BVALID_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic BVALID_param

    );
    export "DPI-C" function axi_initialise_BVALID_from_CY;

    import "DPI-C" context function void axi_set_BRESP_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [1:0] BRESP_param
    );
    import "DPI-C" context function void axi_propagate_BRESP_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BRESP_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [1:0] BRESP_param

    );
    export "DPI-C" function axi_initialise_BRESP_from_CY;

    import "DPI-C" context function void axi_set_BID_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input logic  BID_param
    );
    import "DPI-C" context function void axi_propagate_BID_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BID_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_BID_from_CY_index1;
    export "DPI-C" function axi_initialise_BID_from_CY;

    import "DPI-C" context function void axi_set_BREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic BREADY_param
    );
    import "DPI-C" context function void axi_propagate_BREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic BREADY_param

    );
    export "DPI-C" function axi_initialise_BREADY_from_CY;

    import "DPI-C" context function void axi_set_BUSER_from_SystemVerilog
    (
        input longint _iface_ref,
        input logic [7:0] BUSER_param
    );
    import "DPI-C" context function void axi_propagate_BUSER_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_BUSER_into_SystemVerilog
    (
        input longint _iface_ref,
        output logic [7:0] BUSER_param

    );
    export "DPI-C" function axi_initialise_BUSER_from_CY;

    import "DPI-C" context function void axi_set_config_write_ctrl_to_data_mintime_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_write_ctrl_to_data_mintime_param
    );
    import "DPI-C" context function void axi_propagate_config_write_ctrl_to_data_mintime_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_write_ctrl_to_data_mintime_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_write_ctrl_to_data_mintime_param

    );
    export "DPI-C" function axi_set_config_write_ctrl_to_data_mintime_from_CY;

    import "DPI-C" context function void axi_set_config_master_write_delay_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_master_write_delay_param
    );
    import "DPI-C" context function void axi_propagate_config_master_write_delay_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_deprecated_config_master_write_delay_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_master_write_delay_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_master_write_delay_param

    );
    export "DPI-C" function axi_set_config_master_write_delay_from_CY;

    import "DPI-C" context function void axi_set_config_enable_all_assertions_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_enable_all_assertions_param
    );
    import "DPI-C" context function void axi_propagate_config_enable_all_assertions_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_enable_all_assertions_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_enable_all_assertions_param

    );
    export "DPI-C" function axi_set_config_enable_all_assertions_from_CY;

    import "DPI-C" context function void axi_set_config_enable_assertion_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param
    );
    import "DPI-C" context function void axi_propagate_config_enable_assertion_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_enable_assertion_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param

    );
    export "DPI-C" function axi_set_config_enable_assertion_from_CY;

    import "DPI-C" context function void axi_set_config_slave_start_addr_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input bit  config_slave_start_addr_param
    );
    import "DPI-C" context function void axi_propagate_config_slave_start_addr_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_deprecated_config_slave_start_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_slave_start_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_config_slave_start_addr_from_CY_index1;

    import "DPI-C" context function void axi_set_config_slave_end_addr_from_SystemVerilog_index1
    (
        input longint _iface_ref,
        input int unsigned _this_dot_1,
        input bit  config_slave_end_addr_param
    );
    import "DPI-C" context function void axi_propagate_config_slave_end_addr_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_deprecated_config_slave_end_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_slave_end_addr_into_SystemVerilog
    (
        input longint _iface_ref
    );
    export "DPI-C" function axi_set_config_slave_end_addr_from_CY_index1;

    import "DPI-C" context function void axi_set_config_support_exclusive_access_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_support_exclusive_access_param
    );
    import "DPI-C" context function void axi_propagate_config_support_exclusive_access_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_support_exclusive_access_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_support_exclusive_access_param

    );
    export "DPI-C" function axi_set_config_support_exclusive_access_from_CY;

    import "DPI-C" context function void axi_set_config_read_data_reordering_depth_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_read_data_reordering_depth_param
    );
    import "DPI-C" context function void axi_propagate_config_read_data_reordering_depth_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_read_data_reordering_depth_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_read_data_reordering_depth_param

    );
    export "DPI-C" function axi_set_config_read_data_reordering_depth_from_CY;

    import "DPI-C" context function void axi_set_config_max_transaction_time_factor_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_transaction_time_factor_param
    );
    import "DPI-C" context function void axi_propagate_config_max_transaction_time_factor_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_transaction_time_factor_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_transaction_time_factor_param

    );
    export "DPI-C" function axi_set_config_max_transaction_time_factor_from_CY;

    import "DPI-C" context function void axi_set_config_timeout_max_data_transfer_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_timeout_max_data_transfer_param
    );
    import "DPI-C" context function void axi_propagate_config_timeout_max_data_transfer_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_timeout_max_data_transfer_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_timeout_max_data_transfer_param

    );
    export "DPI-C" function axi_set_config_timeout_max_data_transfer_from_CY;

    import "DPI-C" context function void axi_set_config_burst_timeout_factor_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_burst_timeout_factor_param
    );
    import "DPI-C" context function void axi_propagate_config_burst_timeout_factor_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_burst_timeout_factor_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_burst_timeout_factor_param

    );
    export "DPI-C" function axi_set_config_burst_timeout_factor_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_AWVALID_assertion_to_AWREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_AWVALID_assertion_to_AWREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_ARVALID_assertion_to_ARREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_ARVALID_assertion_to_ARREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_RVALID_assertion_to_RREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_RVALID_assertion_to_RREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_RVALID_assertion_to_RREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_RVALID_assertion_to_RREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_BVALID_assertion_to_BREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_BVALID_assertion_to_BREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_BVALID_assertion_to_BREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_BVALID_assertion_to_BREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_CY;

    import "DPI-C" context function void axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog
    (
        input longint _iface_ref,
        input int unsigned config_max_latency_WVALID_assertion_to_WREADY_param
    );
    import "DPI-C" context function void axi_propagate_config_max_latency_WVALID_assertion_to_WREADY_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_latency_WVALID_assertion_to_WREADY_into_SystemVerilog
    (
        input longint _iface_ref,
        output int unsigned config_max_latency_WVALID_assertion_to_WREADY_param

    );
    export "DPI-C" function axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_CY;

    import "DPI-C" context function void axi_set_config_master_error_position_from_SystemVerilog
    (
        input longint _iface_ref,
        input axi_error_e config_master_error_position_param
    );
    import "DPI-C" context function void axi_propagate_config_master_error_position_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_deprecated_config_master_error_position_into_SystemVerilog
    (
        input longint _iface_ref
    );
    import "DPI-C" context function void axi_get_config_master_error_position_into_SystemVerilog
    (
        input longint _iface_ref,
        output axi_error_e config_master_error_position_param

    );
    export "DPI-C" function axi_set_config_master_error_position_from_CY;

    import "DPI-C" context function void axi_set_config_setup_time_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_setup_time_param
    );
    import "DPI-C" context function void axi_propagate_config_setup_time_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_setup_time_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_setup_time_param

    );
    export "DPI-C" function axi_set_config_setup_time_from_CY;

    import "DPI-C" context function void axi_set_config_hold_time_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_hold_time_param
    );
    import "DPI-C" context function void axi_propagate_config_hold_time_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_hold_time_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_hold_time_param

    );
    export "DPI-C" function axi_set_config_hold_time_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_wr_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_wr_param
    );
    import "DPI-C" context function void axi_propagate_config_max_outstanding_wr_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_outstanding_wr_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_wr_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_wr_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_rd_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_rd_param
    );
    import "DPI-C" context function void axi_propagate_config_max_outstanding_rd_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_outstanding_rd_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_rd_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_rd_from_CY;

    import "DPI-C" context function void axi_set_config_max_outstanding_rw_from_SystemVerilog
    (
        input longint _iface_ref,
        input int config_max_outstanding_rw_param
    );
    import "DPI-C" context function void axi_propagate_config_max_outstanding_rw_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_max_outstanding_rw_into_SystemVerilog
    (
        input longint _iface_ref,
        output int config_max_outstanding_rw_param

    );
    export "DPI-C" function axi_set_config_max_outstanding_rw_from_CY;

    import "DPI-C" context function void axi_set_config_is_issuing_from_SystemVerilog
    (
        input longint _iface_ref,
        input bit config_is_issuing_param
    );
    import "DPI-C" context function void axi_propagate_config_is_issuing_from_SystemVerilog
    (
        input longint _iface_ref    );
    import "DPI-C" context function void axi_get_config_is_issuing_into_SystemVerilog
    (
        input longint _iface_ref,
        output bit config_is_issuing_param

    );
    export "DPI-C" function axi_set_config_is_issuing_from_CY;

    function void axi_initialise_ACLK_from_CY();
        internal_ACLK = 'z;
        m_ACLK = 'z;
    endfunction

    function void axi_initialise_ARESETn_from_CY();
        internal_ARESETn = 'z;
        m_ARESETn = 'z;
    endfunction

    function void axi_initialise_AWVALID_from_CY();
        internal_AWVALID = 'z;
        m_AWVALID = 'z;
    endfunction

    function void axi_set_AWADDR_from_CY_index1( int _this_dot_1, logic  AWADDR_param );
        internal_AWADDR[_this_dot_1] = AWADDR_param;
    endfunction

    function void axi_initialise_AWADDR_from_CY();
        internal_AWADDR = 'z;
        m_AWADDR = 'z;
    endfunction

    function void axi_initialise_AWLEN_from_CY();
        internal_AWLEN = 'z;
        m_AWLEN = 'z;
    endfunction

    function void axi_initialise_AWSIZE_from_CY();
        internal_AWSIZE = 'z;
        m_AWSIZE = 'z;
    endfunction

    function void axi_initialise_AWBURST_from_CY();
        internal_AWBURST = 'z;
        m_AWBURST = 'z;
    endfunction

    function void axi_initialise_AWLOCK_from_CY();
        internal_AWLOCK = 'z;
        m_AWLOCK = 'z;
    endfunction

    function void axi_initialise_AWCACHE_from_CY();
        internal_AWCACHE = 'z;
        m_AWCACHE = 'z;
    endfunction

    function void axi_initialise_AWPROT_from_CY();
        internal_AWPROT = 'z;
        m_AWPROT = 'z;
    endfunction

    function void axi_set_AWID_from_CY_index1( int _this_dot_1, logic  AWID_param );
        internal_AWID[_this_dot_1] = AWID_param;
    endfunction

    function void axi_initialise_AWID_from_CY();
        internal_AWID = 'z;
        m_AWID = 'z;
    endfunction

    function void axi_initialise_AWREADY_from_CY();
        internal_AWREADY = 'z;
        m_AWREADY = 'z;
    endfunction

    function void axi_initialise_AWUSER_from_CY();
        internal_AWUSER = 'z;
        m_AWUSER = 'z;
    endfunction

    function void axi_initialise_ARVALID_from_CY();
        internal_ARVALID = 'z;
        m_ARVALID = 'z;
    endfunction

    function void axi_set_ARADDR_from_CY_index1( int _this_dot_1, logic  ARADDR_param );
        internal_ARADDR[_this_dot_1] = ARADDR_param;
    endfunction

    function void axi_initialise_ARADDR_from_CY();
        internal_ARADDR = 'z;
        m_ARADDR = 'z;
    endfunction

    function void axi_initialise_ARLEN_from_CY();
        internal_ARLEN = 'z;
        m_ARLEN = 'z;
    endfunction

    function void axi_initialise_ARSIZE_from_CY();
        internal_ARSIZE = 'z;
        m_ARSIZE = 'z;
    endfunction

    function void axi_initialise_ARBURST_from_CY();
        internal_ARBURST = 'z;
        m_ARBURST = 'z;
    endfunction

    function void axi_initialise_ARLOCK_from_CY();
        internal_ARLOCK = 'z;
        m_ARLOCK = 'z;
    endfunction

    function void axi_initialise_ARCACHE_from_CY();
        internal_ARCACHE = 'z;
        m_ARCACHE = 'z;
    endfunction

    function void axi_initialise_ARPROT_from_CY();
        internal_ARPROT = 'z;
        m_ARPROT = 'z;
    endfunction

    function void axi_set_ARID_from_CY_index1( int _this_dot_1, logic  ARID_param );
        internal_ARID[_this_dot_1] = ARID_param;
    endfunction

    function void axi_initialise_ARID_from_CY();
        internal_ARID = 'z;
        m_ARID = 'z;
    endfunction

    function void axi_initialise_ARREADY_from_CY();
        internal_ARREADY = 'z;
        m_ARREADY = 'z;
    endfunction

    function void axi_initialise_ARUSER_from_CY();
        internal_ARUSER = 'z;
        m_ARUSER = 'z;
    endfunction

    function void axi_initialise_RVALID_from_CY();
        internal_RVALID = 'z;
        m_RVALID = 'z;
    endfunction

    function void axi_initialise_RLAST_from_CY();
        internal_RLAST = 'z;
        m_RLAST = 'z;
    endfunction

    function void axi_set_RDATA_from_CY_index1( int _this_dot_1, logic  RDATA_param );
        internal_RDATA[_this_dot_1] = RDATA_param;
    endfunction

    function void axi_initialise_RDATA_from_CY();
        internal_RDATA = 'z;
        m_RDATA = 'z;
    endfunction

    function void axi_initialise_RRESP_from_CY();
        internal_RRESP = 'z;
        m_RRESP = 'z;
    endfunction

    function void axi_set_RID_from_CY_index1( int _this_dot_1, logic  RID_param );
        internal_RID[_this_dot_1] = RID_param;
    endfunction

    function void axi_initialise_RID_from_CY();
        internal_RID = 'z;
        m_RID = 'z;
    endfunction

    function void axi_initialise_RREADY_from_CY();
        internal_RREADY = 'z;
        m_RREADY = 'z;
    endfunction

    function void axi_initialise_RUSER_from_CY();
        internal_RUSER = 'z;
        m_RUSER = 'z;
    endfunction

    function void axi_initialise_WVALID_from_CY();
        internal_WVALID = 'z;
        m_WVALID = 'z;
    endfunction

    function void axi_initialise_WLAST_from_CY();
        internal_WLAST = 'z;
        m_WLAST = 'z;
    endfunction

    function void axi_set_WDATA_from_CY_index1( int _this_dot_1, logic  WDATA_param );
        internal_WDATA[_this_dot_1] = WDATA_param;
    endfunction

    function void axi_initialise_WDATA_from_CY();
        internal_WDATA = 'z;
        m_WDATA = 'z;
    endfunction

    function void axi_set_WSTRB_from_CY_index1( int _this_dot_1, logic  WSTRB_param );
        internal_WSTRB[_this_dot_1] = WSTRB_param;
    endfunction

    function void axi_initialise_WSTRB_from_CY();
        internal_WSTRB = 'z;
        m_WSTRB = 'z;
    endfunction

    function void axi_set_WID_from_CY_index1( int _this_dot_1, logic  WID_param );
        internal_WID[_this_dot_1] = WID_param;
    endfunction

    function void axi_initialise_WID_from_CY();
        internal_WID = 'z;
        m_WID = 'z;
    endfunction

    function void axi_initialise_WREADY_from_CY();
        internal_WREADY = 'z;
        m_WREADY = 'z;
    endfunction

    function void axi_initialise_WUSER_from_CY();
        internal_WUSER = 'z;
        m_WUSER = 'z;
    endfunction

    function void axi_initialise_BVALID_from_CY();
        internal_BVALID = 'z;
        m_BVALID = 'z;
    endfunction

    function void axi_initialise_BRESP_from_CY();
        internal_BRESP = 'z;
        m_BRESP = 'z;
    endfunction

    function void axi_set_BID_from_CY_index1( int _this_dot_1, logic  BID_param );
        internal_BID[_this_dot_1] = BID_param;
    endfunction

    function void axi_initialise_BID_from_CY();
        internal_BID = 'z;
        m_BID = 'z;
    endfunction

    function void axi_initialise_BREADY_from_CY();
        internal_BREADY = 'z;
        m_BREADY = 'z;
    endfunction

    function void axi_initialise_BUSER_from_CY();
        internal_BUSER = 'z;
        m_BUSER = 'z;
    endfunction

    function void axi_set_config_write_ctrl_to_data_mintime_from_CY( int unsigned config_write_ctrl_to_data_mintime_param );
        config_write_ctrl_to_data_mintime = config_write_ctrl_to_data_mintime_param;
    endfunction

    function void axi_set_config_master_write_delay_from_CY( bit config_master_write_delay_param );
        config_master_write_delay = config_master_write_delay_param;
    endfunction

    function void axi_set_config_enable_all_assertions_from_CY( bit config_enable_all_assertions_param );
        config_enable_all_assertions = config_enable_all_assertions_param;
    endfunction

    function void axi_set_config_enable_assertion_from_CY( bit [(((AXI_COMBINED_ACCEPTANCE_CAPABILITY_VIOLATION + 1)) - 1):0]  config_enable_assertion_param );
        config_enable_assertion = config_enable_assertion_param;
    endfunction

    function void axi_set_config_slave_start_addr_from_CY_index1( int _this_dot_1, bit  config_slave_start_addr_param );
        config_slave_start_addr[_this_dot_1] = config_slave_start_addr_param;
    endfunction

    function void axi_set_config_slave_end_addr_from_CY_index1( int _this_dot_1, bit  config_slave_end_addr_param );
        config_slave_end_addr[_this_dot_1] = config_slave_end_addr_param;
    endfunction

    function void axi_set_config_support_exclusive_access_from_CY( bit config_support_exclusive_access_param );
        config_support_exclusive_access = config_support_exclusive_access_param;
    endfunction

    function void axi_set_config_read_data_reordering_depth_from_CY( int unsigned config_read_data_reordering_depth_param );
        config_read_data_reordering_depth = config_read_data_reordering_depth_param;
    endfunction

    function void axi_set_config_max_transaction_time_factor_from_CY( int unsigned config_max_transaction_time_factor_param );
        config_max_transaction_time_factor = config_max_transaction_time_factor_param;
    endfunction

    function void axi_set_config_timeout_max_data_transfer_from_CY( int config_timeout_max_data_transfer_param );
        config_timeout_max_data_transfer = config_timeout_max_data_transfer_param;
    endfunction

    function void axi_set_config_burst_timeout_factor_from_CY( int unsigned config_burst_timeout_factor_param );
        config_burst_timeout_factor = config_burst_timeout_factor_param;
    endfunction

    function void axi_set_config_max_latency_AWVALID_assertion_to_AWREADY_from_CY( int unsigned config_max_latency_AWVALID_assertion_to_AWREADY_param );
        config_max_latency_AWVALID_assertion_to_AWREADY = config_max_latency_AWVALID_assertion_to_AWREADY_param;
    endfunction

    function void axi_set_config_max_latency_ARVALID_assertion_to_ARREADY_from_CY( int unsigned config_max_latency_ARVALID_assertion_to_ARREADY_param );
        config_max_latency_ARVALID_assertion_to_ARREADY = config_max_latency_ARVALID_assertion_to_ARREADY_param;
    endfunction

    function void axi_set_config_max_latency_RVALID_assertion_to_RREADY_from_CY( int unsigned config_max_latency_RVALID_assertion_to_RREADY_param );
        config_max_latency_RVALID_assertion_to_RREADY = config_max_latency_RVALID_assertion_to_RREADY_param;
    endfunction

    function void axi_set_config_max_latency_BVALID_assertion_to_BREADY_from_CY( int unsigned config_max_latency_BVALID_assertion_to_BREADY_param );
        config_max_latency_BVALID_assertion_to_BREADY = config_max_latency_BVALID_assertion_to_BREADY_param;
    endfunction

    function void axi_set_config_max_latency_WVALID_assertion_to_WREADY_from_CY( int unsigned config_max_latency_WVALID_assertion_to_WREADY_param );
        config_max_latency_WVALID_assertion_to_WREADY = config_max_latency_WVALID_assertion_to_WREADY_param;
    endfunction

    function void axi_set_config_master_error_position_from_CY( axi_error_e config_master_error_position_param );
        config_master_error_position = config_master_error_position_param;
    endfunction

    function void axi_set_config_setup_time_from_CY( int config_setup_time_param );
        config_setup_time = config_setup_time_param;
    endfunction

    function void axi_set_config_hold_time_from_CY( int config_hold_time_param );
        config_hold_time = config_hold_time_param;
    endfunction

    function void axi_set_config_max_outstanding_wr_from_CY( int config_max_outstanding_wr_param );
        config_max_outstanding_wr = config_max_outstanding_wr_param;
    endfunction

    function void axi_set_config_max_outstanding_rd_from_CY( int config_max_outstanding_rd_param );
        config_max_outstanding_rd = config_max_outstanding_rd_param;
    endfunction

    function void axi_set_config_max_outstanding_rw_from_CY( int config_max_outstanding_rw_param );
        config_max_outstanding_rw = config_max_outstanding_rw_param;
    endfunction

    function void axi_set_config_is_issuing_from_CY( bit config_is_issuing_param );
        config_is_issuing = config_is_issuing_param;
    endfunction



    //--------------------------------------------------------------------------
    //
    // Group:- TLM Interface Support
    //
    //--------------------------------------------------------------------------
    export "DPI-C" axi_get_temp_static_rw_transaction_addr = function axi_get_temp_static_rw_transaction_addr;
    export "DPI-C" axi_set_temp_static_rw_transaction_addr = function axi_set_temp_static_rw_transaction_addr;
    export "DPI-C" axi_get_temp_static_rw_transaction_id = function axi_get_temp_static_rw_transaction_id;
    export "DPI-C" axi_set_temp_static_rw_transaction_id = function axi_set_temp_static_rw_transaction_id;
    export "DPI-C" axi_get_temp_static_rw_transaction_data_words = function axi_get_temp_static_rw_transaction_data_words;
    export "DPI-C" axi_set_temp_static_rw_transaction_data_words = function axi_set_temp_static_rw_transaction_data_words;
    export "DPI-C" axi_get_temp_static_rw_transaction_write_strobes = function axi_get_temp_static_rw_transaction_write_strobes;
    export "DPI-C" axi_set_temp_static_rw_transaction_write_strobes = function axi_set_temp_static_rw_transaction_write_strobes;
    export "DPI-C" axi_get_temp_static_rw_transaction_resp = function axi_get_temp_static_rw_transaction_resp;
    export "DPI-C" axi_set_temp_static_rw_transaction_resp = function axi_set_temp_static_rw_transaction_resp;
    export "DPI-C" axi_get_temp_static_rw_transaction_data_user = function axi_get_temp_static_rw_transaction_data_user;
    export "DPI-C" axi_set_temp_static_rw_transaction_data_user = function axi_set_temp_static_rw_transaction_data_user;
    export "DPI-C" axi_get_temp_static_rw_transaction_write_data_beats_delay = function axi_get_temp_static_rw_transaction_write_data_beats_delay;
    export "DPI-C" axi_set_temp_static_rw_transaction_write_data_beats_delay = function axi_set_temp_static_rw_transaction_write_data_beats_delay;
    export "DPI-C" axi_get_temp_static_rw_transaction_data_valid_delay = function axi_get_temp_static_rw_transaction_data_valid_delay;
    export "DPI-C" axi_set_temp_static_rw_transaction_data_valid_delay = function axi_set_temp_static_rw_transaction_data_valid_delay;
    export "DPI-C" axi_get_temp_static_rw_transaction_data_ready_delay = function axi_get_temp_static_rw_transaction_data_ready_delay;
    export "DPI-C" axi_set_temp_static_rw_transaction_data_ready_delay = function axi_set_temp_static_rw_transaction_data_ready_delay;
    import "DPI-C" context axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog =
    task axi_rw_transaction_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [3:0] burst_length,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] addr_user,
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout axi_rw_e read_or_write,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_valid_delay,
        inout int data_valid_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_response_valid_delay,
        inout int address_ready_delay,
        inout int data_ready_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_response_ready_delay,
        inout bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_rw_transaction_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((4) - 1):0] burst_length,
        inout bit [((8) - 1):0] addr_user,
        inout bit [((8) - 1):0] resp_user,
        inout axi_rw_e read_or_write,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int address_valid_delay,
        inout int write_response_valid_delay,
        inout int address_ready_delay,
        inout int write_response_ready_delay,
        inout bit write_data_with_address,
        input int _unit_id
    );
    import "DPI-C" context axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog =
    task axi_rw_transaction_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_valid_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_ready_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_rw_transaction_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((4) - 1):0] burst_length,
        output bit [((8) - 1):0] addr_user,
        output bit [((8) - 1):0] resp_user,
        output axi_rw_e read_or_write,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        output int address_valid_delay,
        output int write_response_valid_delay,
        output int address_ready_delay,
        output int write_response_ready_delay,
        output bit write_data_with_address,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_AXI_read_addr = function axi_get_temp_static_AXI_read_addr;
    export "DPI-C" axi_set_temp_static_AXI_read_addr = function axi_set_temp_static_AXI_read_addr;
    export "DPI-C" axi_get_temp_static_AXI_read_id = function axi_get_temp_static_AXI_read_id;
    export "DPI-C" axi_set_temp_static_AXI_read_id = function axi_set_temp_static_AXI_read_id;
    export "DPI-C" axi_get_temp_static_AXI_read_data_words = function axi_get_temp_static_AXI_read_data_words;
    export "DPI-C" axi_set_temp_static_AXI_read_data_words = function axi_set_temp_static_AXI_read_data_words;
    export "DPI-C" axi_get_temp_static_AXI_read_resp = function axi_get_temp_static_AXI_read_resp;
    export "DPI-C" axi_set_temp_static_AXI_read_resp = function axi_set_temp_static_AXI_read_resp;
    export "DPI-C" axi_get_temp_static_AXI_read_data_user = function axi_get_temp_static_AXI_read_data_user;
    export "DPI-C" axi_set_temp_static_AXI_read_data_user = function axi_set_temp_static_AXI_read_data_user;
    export "DPI-C" axi_get_temp_static_AXI_read_data_start_time = function axi_get_temp_static_AXI_read_data_start_time;
    export "DPI-C" axi_set_temp_static_AXI_read_data_start_time = function axi_set_temp_static_AXI_read_data_start_time;
    export "DPI-C" axi_get_temp_static_AXI_read_data_end_time = function axi_get_temp_static_AXI_read_data_end_time;
    export "DPI-C" axi_set_temp_static_AXI_read_data_end_time = function axi_set_temp_static_AXI_read_data_end_time;
    import "DPI-C" context axi_AXI_read_ActivatesActivatingActivate_SystemVerilog =
    task axi_AXI_read_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [3:0] burst_length,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] addr_user,
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_to_data_latency,
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_AXI_read_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((4) - 1):0] burst_length,
        inout bit [((8) - 1):0] addr_user,
        inout int address_to_data_latency,
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_read_ReceivedReceivingReceive_SystemVerilog =
    task axi_AXI_read_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_AXI_read_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((4) - 1):0] burst_length,
        output bit [((8) - 1):0] addr_user,
        output int address_to_data_latency,
        output longint addr_start_time,
        output longint addr_end_time,
        output int address_valid_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_AXI_write_addr = function axi_get_temp_static_AXI_write_addr;
    export "DPI-C" axi_set_temp_static_AXI_write_addr = function axi_set_temp_static_AXI_write_addr;
    export "DPI-C" axi_get_temp_static_AXI_write_id = function axi_get_temp_static_AXI_write_id;
    export "DPI-C" axi_set_temp_static_AXI_write_id = function axi_set_temp_static_AXI_write_id;
    export "DPI-C" axi_get_temp_static_AXI_write_data_words = function axi_get_temp_static_AXI_write_data_words;
    export "DPI-C" axi_set_temp_static_AXI_write_data_words = function axi_set_temp_static_AXI_write_data_words;
    export "DPI-C" axi_get_temp_static_AXI_write_write_strobes = function axi_get_temp_static_AXI_write_write_strobes;
    export "DPI-C" axi_set_temp_static_AXI_write_write_strobes = function axi_set_temp_static_AXI_write_write_strobes;
    export "DPI-C" axi_get_temp_static_AXI_write_data_user = function axi_get_temp_static_AXI_write_data_user;
    export "DPI-C" axi_set_temp_static_AXI_write_data_user = function axi_set_temp_static_AXI_write_data_user;
    export "DPI-C" axi_get_temp_static_AXI_write_write_data_beats_delay = function axi_get_temp_static_AXI_write_write_data_beats_delay;
    export "DPI-C" axi_set_temp_static_AXI_write_write_data_beats_delay = function axi_set_temp_static_AXI_write_write_data_beats_delay;
    export "DPI-C" axi_get_temp_static_AXI_write_data_start_time = function axi_get_temp_static_AXI_write_data_start_time;
    export "DPI-C" axi_set_temp_static_AXI_write_data_start_time = function axi_set_temp_static_AXI_write_data_start_time;
    export "DPI-C" axi_get_temp_static_AXI_write_data_end_time = function axi_get_temp_static_AXI_write_data_end_time;
    export "DPI-C" axi_set_temp_static_AXI_write_data_end_time = function axi_set_temp_static_AXI_write_data_end_time;
    import "DPI-C" context axi_AXI_write_ActivatesActivatingActivate_SystemVerilog =
    task axi_AXI_write_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [3:0] burst_length,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout axi_response_e resp,
        inout bit [7:0] addr_user,
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint wr_resp_start_time,
        inout longint wr_resp_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_AXI_write_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout axi_size_e size,
        inout axi_burst_e burst,
        inout axi_lock_e lock,
        inout axi_cache_e cache,
        inout axi_prot_e prot,
        inout bit [((4) - 1):0] burst_length,
        inout axi_response_e resp,
        inout bit [((8) - 1):0] addr_user,
        inout bit [((8) - 1):0] resp_user,
        inout int address_to_data_latency,
        inout int data_to_response_latency,
        inout int write_address_to_data_delay,
        inout int write_data_to_address_delay,
        inout longint addr_start_time,
        inout longint addr_end_time,
        inout longint wr_resp_start_time,
        inout longint wr_resp_end_time,
        inout int address_valid_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_AXI_write_ReceivedReceivingReceive_SystemVerilog =
    task axi_AXI_write_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_AXI_write_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((4) - 1):0] burst_length,
        output axi_response_e resp,
        output bit [((8) - 1):0] addr_user,
        output bit [((8) - 1):0] resp_user,
        output int address_to_data_latency,
        output int data_to_response_latency,
        output int write_address_to_data_delay,
        output int write_data_to_address_delay,
        output longint addr_start_time,
        output longint addr_end_time,
        output longint wr_resp_start_time,
        output longint wr_resp_end_time,
        output int address_valid_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_data_resp_data_words = function axi_get_temp_static_data_resp_data_words;
    export "DPI-C" axi_set_temp_static_data_resp_data_words = function axi_set_temp_static_data_resp_data_words;
    export "DPI-C" axi_get_temp_static_data_resp_write_strobes = function axi_get_temp_static_data_resp_write_strobes;
    export "DPI-C" axi_set_temp_static_data_resp_write_strobes = function axi_set_temp_static_data_resp_write_strobes;
    export "DPI-C" axi_get_temp_static_data_resp_id = function axi_get_temp_static_data_resp_id;
    export "DPI-C" axi_set_temp_static_data_resp_id = function axi_set_temp_static_data_resp_id;
    export "DPI-C" axi_get_temp_static_data_resp_data_user = function axi_get_temp_static_data_resp_data_user;
    export "DPI-C" axi_set_temp_static_data_resp_data_user = function axi_set_temp_static_data_resp_data_user;
    export "DPI-C" axi_get_temp_static_data_resp_write_data_beats_delay = function axi_get_temp_static_data_resp_write_data_beats_delay;
    export "DPI-C" axi_set_temp_static_data_resp_write_data_beats_delay = function axi_set_temp_static_data_resp_write_data_beats_delay;
    export "DPI-C" axi_get_temp_static_data_resp_data_beat_start_time = function axi_get_temp_static_data_resp_data_beat_start_time;
    export "DPI-C" axi_set_temp_static_data_resp_data_beat_start_time = function axi_set_temp_static_data_resp_data_beat_start_time;
    export "DPI-C" axi_get_temp_static_data_resp_data_beat_end_time = function axi_get_temp_static_data_resp_data_beat_end_time;
    export "DPI-C" axi_set_temp_static_data_resp_data_beat_end_time = function axi_set_temp_static_data_resp_data_beat_end_time;
    import "DPI-C" context axi_data_resp_ActivatesActivatingActivate_SystemVerilog =
    task axi_data_resp_ActivatesActivatingActivate_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int burst_length,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout axi_response_e resp,
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout bit [7:0] resp_user,
        inout longint data_start,
        inout longint data_end,
        inout longint response_start,
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog =
    task axi_data_resp_ActivatesActivatingActivate_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        inout int burst_length,
        inout axi_response_e resp,
        inout bit [((8) - 1):0] resp_user,
        inout longint data_start,
        inout longint data_end,
        inout longint response_start,
        inout longint response_end_time,
        input int _unit_id
    );
    import "DPI-C" context axi_data_resp_ReceivedReceivingReceive_SystemVerilog =
    task axi_data_resp_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_beat_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_data_resp_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output int burst_length,
        output axi_response_e resp,
        output bit [((8) - 1):0] resp_user,
        output longint data_start,
        output longint data_end,
        output longint response_start,
        output longint response_end_time,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_data_burst_data_words = function axi_get_temp_static_read_data_burst_data_words;
    export "DPI-C" axi_set_temp_static_read_data_burst_data_words = function axi_set_temp_static_read_data_burst_data_words;
    export "DPI-C" axi_get_temp_static_read_data_burst_resp = function axi_get_temp_static_read_data_burst_resp;
    export "DPI-C" axi_set_temp_static_read_data_burst_resp = function axi_set_temp_static_read_data_burst_resp;
    export "DPI-C" axi_get_temp_static_read_data_burst_id = function axi_get_temp_static_read_data_burst_id;
    export "DPI-C" axi_set_temp_static_read_data_burst_id = function axi_set_temp_static_read_data_burst_id;
    export "DPI-C" axi_get_temp_static_read_data_burst_data_user = function axi_get_temp_static_read_data_burst_data_user;
    export "DPI-C" axi_set_temp_static_read_data_burst_data_user = function axi_set_temp_static_read_data_burst_data_user;
    export "DPI-C" axi_get_temp_static_read_data_burst_data_start_time = function axi_get_temp_static_read_data_burst_data_start_time;
    export "DPI-C" axi_set_temp_static_read_data_burst_data_start_time = function axi_set_temp_static_read_data_burst_data_start_time;
    export "DPI-C" axi_get_temp_static_read_data_burst_data_end_time = function axi_get_temp_static_read_data_burst_data_end_time;
    export "DPI-C" axi_set_temp_static_read_data_burst_data_end_time = function axi_set_temp_static_read_data_burst_data_end_time;
    import "DPI-C" context axi_read_data_burst_SendSendingSent_SystemVerilog =
    task axi_read_data_burst_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_data_burst_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int resp_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_data_burst_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_data_burst_data_words = function axi_get_temp_static_write_data_burst_data_words;
    export "DPI-C" axi_set_temp_static_write_data_burst_data_words = function axi_set_temp_static_write_data_burst_data_words;
    export "DPI-C" axi_get_temp_static_write_data_burst_write_strobes = function axi_get_temp_static_write_data_burst_write_strobes;
    export "DPI-C" axi_set_temp_static_write_data_burst_write_strobes = function axi_set_temp_static_write_data_burst_write_strobes;
    export "DPI-C" axi_get_temp_static_write_data_burst_id = function axi_get_temp_static_write_data_burst_id;
    export "DPI-C" axi_set_temp_static_write_data_burst_id = function axi_set_temp_static_write_data_burst_id;
    export "DPI-C" axi_get_temp_static_write_data_burst_data_user = function axi_get_temp_static_write_data_burst_data_user;
    export "DPI-C" axi_set_temp_static_write_data_burst_data_user = function axi_set_temp_static_write_data_burst_data_user;
    export "DPI-C" axi_get_temp_static_write_data_burst_write_data_beats_delay = function axi_get_temp_static_write_data_burst_write_data_beats_delay;
    export "DPI-C" axi_set_temp_static_write_data_burst_write_data_beats_delay = function axi_set_temp_static_write_data_burst_write_data_beats_delay;
    export "DPI-C" axi_get_temp_static_write_data_burst_data_start_time = function axi_get_temp_static_write_data_burst_data_start_time;
    export "DPI-C" axi_set_temp_static_write_data_burst_data_start_time = function axi_set_temp_static_write_data_burst_data_start_time;
    export "DPI-C" axi_get_temp_static_write_data_burst_data_end_time = function axi_get_temp_static_write_data_burst_data_end_time;
    export "DPI-C" axi_set_temp_static_write_data_burst_data_end_time = function axi_set_temp_static_write_data_burst_data_end_time;
    import "DPI-C" context axi_write_data_burst_SendSendingSent_SystemVerilog =
    task axi_write_data_burst_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int burst_length,
        input int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id
    );
    import "DPI-C" context axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_data_burst_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        inout int data_words_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_strobes_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_user_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int write_data_beats_delay_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_start_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        inout int data_end_time_DIMS0, // Array to pass in and/or out the unsized dims of param
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_data_burst_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output int burst_length,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_addr_channel_phase_addr = function axi_get_temp_static_read_addr_channel_phase_addr;
    export "DPI-C" axi_set_temp_static_read_addr_channel_phase_addr = function axi_set_temp_static_read_addr_channel_phase_addr;
    export "DPI-C" axi_get_temp_static_read_addr_channel_phase_id = function axi_get_temp_static_read_addr_channel_phase_id;
    export "DPI-C" axi_set_temp_static_read_addr_channel_phase_id = function axi_set_temp_static_read_addr_channel_phase_id;
    import "DPI-C" context axi_read_addr_channel_phase_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((8) - 1):0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_channel_phase_data = function axi_get_temp_static_read_channel_phase_data;
    export "DPI-C" axi_set_temp_static_read_channel_phase_data = function axi_set_temp_static_read_channel_phase_data;
    export "DPI-C" axi_get_temp_static_read_channel_phase_id = function axi_get_temp_static_read_channel_phase_id;
    export "DPI-C" axi_set_temp_static_read_channel_phase_id = function axi_set_temp_static_read_channel_phase_id;
    import "DPI-C" context axi_read_channel_phase_SendSendingSent_SystemVerilog =
    task axi_read_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input axi_response_e resp,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output axi_response_e resp,
        output bit [((8) - 1):0] data_user,
        output int data_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_addr_channel_phase_addr = function axi_get_temp_static_write_addr_channel_phase_addr;
    export "DPI-C" axi_set_temp_static_write_addr_channel_phase_addr = function axi_set_temp_static_write_addr_channel_phase_addr;
    export "DPI-C" axi_get_temp_static_write_addr_channel_phase_id = function axi_get_temp_static_write_addr_channel_phase_id;
    export "DPI-C" axi_set_temp_static_write_addr_channel_phase_id = function axi_set_temp_static_write_addr_channel_phase_id;
    import "DPI-C" context axi_write_addr_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [7:0] addr_user,
        input int address_valid_delay,
        input int address_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_addr_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((8) - 1):0] addr_user,
        output int address_valid_delay,
        output int address_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_channel_phase_data = function axi_get_temp_static_write_channel_phase_data;
    export "DPI-C" axi_set_temp_static_write_channel_phase_data = function axi_set_temp_static_write_channel_phase_data;
    export "DPI-C" axi_get_temp_static_write_channel_phase_write_strobes = function axi_get_temp_static_write_channel_phase_write_strobes;
    export "DPI-C" axi_set_temp_static_write_channel_phase_write_strobes = function axi_set_temp_static_write_channel_phase_write_strobes;
    export "DPI-C" axi_get_temp_static_write_channel_phase_id = function axi_get_temp_static_write_channel_phase_id;
    export "DPI-C" axi_set_temp_static_write_channel_phase_id = function axi_set_temp_static_write_channel_phase_id;
    import "DPI-C" context axi_write_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [7:0] data_user,
        input int data_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output bit [((8) - 1):0] data_user,
        output int data_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_resp_channel_phase_id = function axi_get_temp_static_write_resp_channel_phase_id;
    export "DPI-C" axi_set_temp_static_write_resp_channel_phase_id = function axi_set_temp_static_write_resp_channel_phase_id;
    import "DPI-C" context axi_write_resp_channel_phase_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_phase_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [7:0] resp_user,
        input int write_response_ready_delay,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_phase_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_phase_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_resp_channel_phase_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_response_e resp,
        output bit [((8) - 1):0] resp_user,
        output int write_response_ready_delay,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_addr_channel_cycle_addr = function axi_get_temp_static_read_addr_channel_cycle_addr;
    export "DPI-C" axi_set_temp_static_read_addr_channel_cycle_addr = function axi_set_temp_static_read_addr_channel_cycle_addr;
    export "DPI-C" axi_get_temp_static_read_addr_channel_cycle_id = function axi_get_temp_static_read_addr_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_read_addr_channel_cycle_id = function axi_set_temp_static_read_addr_channel_cycle_id;
    import "DPI-C" context axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((8) - 1):0] addr_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_addr_channel_ready_SendSendingSent_SystemVerilog =
    task axi_read_addr_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_read_channel_cycle_data = function axi_get_temp_static_read_channel_cycle_data;
    export "DPI-C" axi_set_temp_static_read_channel_cycle_data = function axi_set_temp_static_read_channel_cycle_data;
    export "DPI-C" axi_get_temp_static_read_channel_cycle_id = function axi_get_temp_static_read_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_read_channel_cycle_id = function axi_set_temp_static_read_channel_cycle_id;
    import "DPI-C" context axi_read_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_read_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input axi_response_e resp,
        input bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_read_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output axi_response_e resp,
        output bit [((8) - 1):0] data_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_read_channel_ready_SendSendingSent_SystemVerilog =
    task axi_read_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_read_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_addr_channel_cycle_addr = function axi_get_temp_static_write_addr_channel_cycle_addr;
    export "DPI-C" axi_set_temp_static_write_addr_channel_cycle_addr = function axi_set_temp_static_write_addr_channel_cycle_addr;
    export "DPI-C" axi_get_temp_static_write_addr_channel_cycle_id = function axi_get_temp_static_write_addr_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_write_addr_channel_cycle_id = function axi_set_temp_static_write_addr_channel_cycle_id;
    import "DPI-C" context axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit [3:0] burst_length,
        input axi_size_e size,
        input axi_burst_e burst,
        input axi_lock_e lock,
        input axi_cache_e cache,
        input axi_prot_e prot,
        input bit [7:0] addr_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_addr_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit [((4) - 1):0] burst_length,
        output axi_size_e size,
        output axi_burst_e burst,
        output axi_lock_e lock,
        output axi_cache_e cache,
        output axi_prot_e prot,
        output bit [((8) - 1):0] addr_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_addr_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_addr_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_addr_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_channel_cycle_data = function axi_get_temp_static_write_channel_cycle_data;
    export "DPI-C" axi_set_temp_static_write_channel_cycle_data = function axi_set_temp_static_write_channel_cycle_data;
    export "DPI-C" axi_get_temp_static_write_channel_cycle_strb = function axi_get_temp_static_write_channel_cycle_strb;
    export "DPI-C" axi_set_temp_static_write_channel_cycle_strb = function axi_set_temp_static_write_channel_cycle_strb;
    export "DPI-C" axi_get_temp_static_write_channel_cycle_id = function axi_get_temp_static_write_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_write_channel_cycle_id = function axi_set_temp_static_write_channel_cycle_id;
    import "DPI-C" context axi_write_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit last,
        input bit [7:0] data_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output bit last,
        output bit [((8) - 1):0] data_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    export "DPI-C" axi_get_temp_static_write_resp_channel_cycle_id = function axi_get_temp_static_write_resp_channel_cycle_id;
    export "DPI-C" axi_set_temp_static_write_resp_channel_cycle_id = function axi_set_temp_static_write_resp_channel_cycle_id;
    import "DPI-C" context axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_cycle_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input axi_response_e resp,
        input bit [7:0] resp_user,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_cycle_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output int _trans_id,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog =
    task axi_write_resp_channel_cycle_ReceivedReceivingReceive_open_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input int _trans_id,
        output axi_response_e resp,
        output bit [((8) - 1):0] resp_user,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_write_resp_channel_ready_SendSendingSent_SystemVerilog =
    task axi_write_resp_channel_ready_SendSendingSent_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        input bit ready,
        input int _unit_id
    );
    import "DPI-C" context axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog =
    task axi_write_resp_channel_ready_ReceivedReceivingReceive_SystemVerilog
    (
        input int _comms_semantic,
        input longint _as_end,
        output bit ready,
        input int _unit_id,
        input bit _using
    );
    import "DPI-C" context axi_end_of_timestep_VPI_SystemVerilog =
    task axi_end_of_timestep_VPI_SystemVerilog();
    import "DPI-C" context axi_fn_rd_txn_valid_lanes = function void fn_rd_txn_valid_lanes_C
    (
    );

    import "DPI-C" context axi_fn_get_wdata_phase_info = function void fn_get_wdata_phase_info_C
    (
        input bit wdata_last,
        inout bit waddr_rcvd,
        output bit [3:0] burst_length,
        output int beat_num
    );

    import "DPI-C" context axi_fn_get_wresp_phase_info = function void fn_get_wresp_phase_info_C
    (
    );

    import "DPI-C" context axi_fn_get_rdata_phase_info = function void fn_get_rdata_phase_info_C
    (
        input bit rdata_last,
        output bit [3:0] burst_length,
        output int beat_num
    );

    import "DPI-C" context axi_fn_get_max_os_per_id = function void fn_get_max_os_per_id_C
    (
        output int max_waddr_os,
        output int max_wdata_os
    );

    import "DPI-C" context axi_get_rw_txns_in_prog = function void get_rw_txns_in_prog_C
    (
        output axi_rw_txn_counts_s txn_counts
    );

    import "DPI-C" context axi_fn_add_addr_map_entry = function void fn_add_addr_map_entry_C
    (
        input string region,
        input longint unsigned size
    );

    import "DPI-C" context axi_fn_add_wr_delay = function void fn_add_wr_delay_C
    (
        input string region,
        input bit [17:0] id,
        input int unsigned addr2data,
        input int data2data_DIMS0
    );

    import "DPI-C" context axi_fn_delete_wr_delay = function void fn_delete_wr_delay_C
    (
        input string region,
        input bit [17:0] id
    );

    import "DPI-C" context axi_fn_set_wr_def_delays = function void fn_set_wr_def_delays_C
    (
        input int unsigned min_addr2data,
        input int min_data2data_DIMS0,
        input int unsigned max_addr2data,
        input int max_data2data_DIMS0
    );

    // Waiter task and control
    reg wait_for_control = 0;

    always @(posedge wait_for_control)
    begin
        disable wait_for;
        wait_for_control = 0;
    end

    export "DPI-C" axi_wait_for = task wait_for;

    task wait_for();
        begin
            wait(0 == 1);
        end
    endtask

    // Drive wires (from Cohesive) 
    assign ACLK = internal_ACLK;
    assign ARESETn = internal_ARESETn;
    assign AWVALID = internal_AWVALID;
    assign AWADDR = internal_AWADDR;
    assign AWLEN = internal_AWLEN;
    assign AWSIZE = internal_AWSIZE;
    assign AWBURST = internal_AWBURST;
    assign AWLOCK = internal_AWLOCK;
    assign AWCACHE = internal_AWCACHE;
    assign AWPROT = internal_AWPROT;
    assign AWID = internal_AWID;
    assign AWREADY = internal_AWREADY;
    assign AWUSER = internal_AWUSER;
    assign ARVALID = internal_ARVALID;
    assign ARADDR = internal_ARADDR;
    assign ARLEN = internal_ARLEN;
    assign ARSIZE = internal_ARSIZE;
    assign ARBURST = internal_ARBURST;
    assign ARLOCK = internal_ARLOCK;
    assign ARCACHE = internal_ARCACHE;
    assign ARPROT = internal_ARPROT;
    assign ARID = internal_ARID;
    assign ARREADY = internal_ARREADY;
    assign ARUSER = internal_ARUSER;
    assign RVALID = internal_RVALID;
    assign RLAST = internal_RLAST;
    assign RDATA = internal_RDATA;
    assign RRESP = internal_RRESP;
    assign RID = internal_RID;
    assign RREADY = internal_RREADY;
    assign RUSER = internal_RUSER;
    assign WVALID = internal_WVALID;
    assign WLAST = internal_WLAST;
    assign WDATA = internal_WDATA;
    assign WSTRB = internal_WSTRB;
    assign WID = internal_WID;
    assign WREADY = internal_WREADY;
    assign WUSER = internal_WUSER;
    assign BVALID = internal_BVALID;
    assign BRESP = internal_BRESP;
    assign BID = internal_BID;
    assign BREADY = internal_BREADY;
    assign BUSER = internal_BUSER;
    // Drive wires (from User) 
    assign ACLK = m_ACLK;
    assign ARESETn = m_ARESETn;
    assign AWVALID = m_AWVALID;
    assign AWADDR = m_AWADDR;
    assign AWLEN = m_AWLEN;
    assign AWSIZE = m_AWSIZE;
    assign AWBURST = m_AWBURST;
    assign AWLOCK = m_AWLOCK;
    assign AWCACHE = m_AWCACHE;
    assign AWPROT = m_AWPROT;
    assign AWID = m_AWID;
    assign AWREADY = m_AWREADY;
    assign AWUSER = m_AWUSER;
    assign ARVALID = m_ARVALID;
    assign ARADDR = m_ARADDR;
    assign ARLEN = m_ARLEN;
    assign ARSIZE = m_ARSIZE;
    assign ARBURST = m_ARBURST;
    assign ARLOCK = m_ARLOCK;
    assign ARCACHE = m_ARCACHE;
    assign ARPROT = m_ARPROT;
    assign ARID = m_ARID;
    assign ARREADY = m_ARREADY;
    assign ARUSER = m_ARUSER;
    assign RVALID = m_RVALID;
    assign RLAST = m_RLAST;
    assign RDATA = m_RDATA;
    assign RRESP = m_RRESP;
    assign RID = m_RID;
    assign RREADY = m_RREADY;
    assign RUSER = m_RUSER;
    assign WVALID = m_WVALID;
    assign WLAST = m_WLAST;
    assign WDATA = m_WDATA;
    assign WSTRB = m_WSTRB;
    assign WID = m_WID;
    assign WREADY = m_WREADY;
    assign WUSER = m_WUSER;
    assign BVALID = m_BVALID;
    assign BRESP = m_BRESP;
    assign BID = m_BID;
    assign BREADY = m_BREADY;
    assign BUSER = m_BUSER;

    reg ACLK_changed = 0;
    reg ARESETn_changed = 0;
    reg AWVALID_changed = 0;
    reg AWADDR_changed = 0;
    reg AWLEN_changed = 0;
    reg AWSIZE_changed = 0;
    reg AWBURST_changed = 0;
    reg AWLOCK_changed = 0;
    reg AWCACHE_changed = 0;
    reg AWPROT_changed = 0;
    reg AWID_changed = 0;
    reg AWREADY_changed = 0;
    reg AWUSER_changed = 0;
    reg ARVALID_changed = 0;
    reg ARADDR_changed = 0;
    reg ARLEN_changed = 0;
    reg ARSIZE_changed = 0;
    reg ARBURST_changed = 0;
    reg ARLOCK_changed = 0;
    reg ARCACHE_changed = 0;
    reg ARPROT_changed = 0;
    reg ARID_changed = 0;
    reg ARREADY_changed = 0;
    reg ARUSER_changed = 0;
    reg RVALID_changed = 0;
    reg RLAST_changed = 0;
    reg RDATA_changed = 0;
    reg RRESP_changed = 0;
    reg RID_changed = 0;
    reg RREADY_changed = 0;
    reg RUSER_changed = 0;
    reg WVALID_changed = 0;
    reg WLAST_changed = 0;
    reg WDATA_changed = 0;
    reg WSTRB_changed = 0;
    reg WID_changed = 0;
    reg WREADY_changed = 0;
    reg WUSER_changed = 0;
    reg BVALID_changed = 0;
    reg BRESP_changed = 0;
    reg BID_changed = 0;
    reg BREADY_changed = 0;
    reg BUSER_changed = 0;
    reg config_write_ctrl_to_data_mintime_changed = 0;
    reg config_master_write_delay_changed = 0;
    reg config_enable_all_assertions_changed = 0;
    reg config_enable_assertion_changed = 0;
    reg config_slave_start_addr_changed = 0;
    reg config_slave_end_addr_changed = 0;
    reg config_support_exclusive_access_changed = 0;
    reg config_read_data_reordering_depth_changed = 0;
    reg config_max_transaction_time_factor_changed = 0;
    reg config_timeout_max_data_transfer_changed = 0;
    reg config_burst_timeout_factor_changed = 0;
    reg config_max_latency_AWVALID_assertion_to_AWREADY_changed = 0;
    reg config_max_latency_ARVALID_assertion_to_ARREADY_changed = 0;
    reg config_max_latency_RVALID_assertion_to_RREADY_changed = 0;
    reg config_max_latency_BVALID_assertion_to_BREADY_changed = 0;
    reg config_max_latency_WVALID_assertion_to_WREADY_changed = 0;
    reg config_master_error_position_changed = 0;
    reg config_setup_time_changed = 0;
    reg config_hold_time_changed = 0;
    reg config_max_outstanding_wr_changed = 0;
    reg config_max_outstanding_rd_changed = 0;
    reg config_max_outstanding_rw_changed = 0;
    reg config_is_issuing_changed = 0;

    reg end_of_timestep_control = 0;

    // Start end_of_timestep timer
    initial
    forever
    begin
        wait_end_of_timestep();
    end


    event non_blocking_end_of_timestep_control;

    export "DPI-C" axi_wait_end_of_timestep = task wait_end_of_timestep;

    task wait_end_of_timestep();
        begin
            @(non_blocking_end_of_timestep_control);
            axi_end_of_timestep_VPI_SystemVerilog();
        end
    endtask

    always @( posedge end_of_timestep_control or posedge _check_t0_values )
    begin
        if ( end_of_timestep_control == 1 )
        begin
            ->> non_blocking_end_of_timestep_control;
            end_of_timestep_control = 0;
        end
    end


    // SV wire change monitors

    function automatic void axi_local_set_ACLK_from_SystemVerilog(  );
            axi_set_ACLK_from_SystemVerilog( _interface_ref, ACLK); // DPI call to imported task
        
        axi_propagate_ACLK_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ACLK or posedge _check_t0_values )
    begin
        axi_local_set_ACLK_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARESETn_from_SystemVerilog(  );
            axi_set_ARESETn_from_SystemVerilog( _interface_ref, ARESETn); // DPI call to imported task
        
        axi_propagate_ARESETn_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARESETn or posedge _check_t0_values )
    begin
        axi_local_set_ARESETn_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWVALID_from_SystemVerilog(  );
            axi_set_AWVALID_from_SystemVerilog( _interface_ref, AWVALID); // DPI call to imported task
        
        axi_propagate_AWVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWVALID or posedge _check_t0_values )
    begin
        axi_local_set_AWVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWADDR_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ADDRESS_WIDTH ); _this_dot_1++)
        begin
            axi_set_AWADDR_from_SystemVerilog_index1( _interface_ref, _this_dot_1,AWADDR[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_AWADDR_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWADDR or posedge _check_t0_values )
    begin
        axi_local_set_AWADDR_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWLEN_from_SystemVerilog(  );
            axi_set_AWLEN_from_SystemVerilog( _interface_ref, AWLEN); // DPI call to imported task
        
        axi_propagate_AWLEN_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWLEN or posedge _check_t0_values )
    begin
        axi_local_set_AWLEN_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWSIZE_from_SystemVerilog(  );
            axi_set_AWSIZE_from_SystemVerilog( _interface_ref, AWSIZE); // DPI call to imported task
        
        axi_propagate_AWSIZE_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWSIZE or posedge _check_t0_values )
    begin
        axi_local_set_AWSIZE_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWBURST_from_SystemVerilog(  );
            axi_set_AWBURST_from_SystemVerilog( _interface_ref, AWBURST); // DPI call to imported task
        
        axi_propagate_AWBURST_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWBURST or posedge _check_t0_values )
    begin
        axi_local_set_AWBURST_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWLOCK_from_SystemVerilog(  );
            axi_set_AWLOCK_from_SystemVerilog( _interface_ref, AWLOCK); // DPI call to imported task
        
        axi_propagate_AWLOCK_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWLOCK or posedge _check_t0_values )
    begin
        axi_local_set_AWLOCK_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWCACHE_from_SystemVerilog(  );
            axi_set_AWCACHE_from_SystemVerilog( _interface_ref, AWCACHE); // DPI call to imported task
        
        axi_propagate_AWCACHE_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWCACHE or posedge _check_t0_values )
    begin
        axi_local_set_AWCACHE_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWPROT_from_SystemVerilog(  );
            axi_set_AWPROT_from_SystemVerilog( _interface_ref, AWPROT); // DPI call to imported task
        
        axi_propagate_AWPROT_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWPROT or posedge _check_t0_values )
    begin
        axi_local_set_AWPROT_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_AWID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,AWID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_AWID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWID or posedge _check_t0_values )
    begin
        axi_local_set_AWID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWREADY_from_SystemVerilog(  );
            axi_set_AWREADY_from_SystemVerilog( _interface_ref, AWREADY); // DPI call to imported task
        
        axi_propagate_AWREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWREADY or posedge _check_t0_values )
    begin
        axi_local_set_AWREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_AWUSER_from_SystemVerilog(  );
            axi_set_AWUSER_from_SystemVerilog( _interface_ref, AWUSER); // DPI call to imported task
        
        axi_propagate_AWUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( AWUSER or posedge _check_t0_values )
    begin
        axi_local_set_AWUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARVALID_from_SystemVerilog(  );
            axi_set_ARVALID_from_SystemVerilog( _interface_ref, ARVALID); // DPI call to imported task
        
        axi_propagate_ARVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARVALID or posedge _check_t0_values )
    begin
        axi_local_set_ARVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARADDR_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ADDRESS_WIDTH ); _this_dot_1++)
        begin
            axi_set_ARADDR_from_SystemVerilog_index1( _interface_ref, _this_dot_1,ARADDR[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_ARADDR_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARADDR or posedge _check_t0_values )
    begin
        axi_local_set_ARADDR_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARLEN_from_SystemVerilog(  );
            axi_set_ARLEN_from_SystemVerilog( _interface_ref, ARLEN); // DPI call to imported task
        
        axi_propagate_ARLEN_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARLEN or posedge _check_t0_values )
    begin
        axi_local_set_ARLEN_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARSIZE_from_SystemVerilog(  );
            axi_set_ARSIZE_from_SystemVerilog( _interface_ref, ARSIZE); // DPI call to imported task
        
        axi_propagate_ARSIZE_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARSIZE or posedge _check_t0_values )
    begin
        axi_local_set_ARSIZE_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARBURST_from_SystemVerilog(  );
            axi_set_ARBURST_from_SystemVerilog( _interface_ref, ARBURST); // DPI call to imported task
        
        axi_propagate_ARBURST_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARBURST or posedge _check_t0_values )
    begin
        axi_local_set_ARBURST_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARLOCK_from_SystemVerilog(  );
            axi_set_ARLOCK_from_SystemVerilog( _interface_ref, ARLOCK); // DPI call to imported task
        
        axi_propagate_ARLOCK_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARLOCK or posedge _check_t0_values )
    begin
        axi_local_set_ARLOCK_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARCACHE_from_SystemVerilog(  );
            axi_set_ARCACHE_from_SystemVerilog( _interface_ref, ARCACHE); // DPI call to imported task
        
        axi_propagate_ARCACHE_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARCACHE or posedge _check_t0_values )
    begin
        axi_local_set_ARCACHE_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARPROT_from_SystemVerilog(  );
            axi_set_ARPROT_from_SystemVerilog( _interface_ref, ARPROT); // DPI call to imported task
        
        axi_propagate_ARPROT_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARPROT or posedge _check_t0_values )
    begin
        axi_local_set_ARPROT_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_ARID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,ARID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_ARID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARID or posedge _check_t0_values )
    begin
        axi_local_set_ARID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARREADY_from_SystemVerilog(  );
            axi_set_ARREADY_from_SystemVerilog( _interface_ref, ARREADY); // DPI call to imported task
        
        axi_propagate_ARREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARREADY or posedge _check_t0_values )
    begin
        axi_local_set_ARREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_ARUSER_from_SystemVerilog(  );
            axi_set_ARUSER_from_SystemVerilog( _interface_ref, ARUSER); // DPI call to imported task
        
        axi_propagate_ARUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( ARUSER or posedge _check_t0_values )
    begin
        axi_local_set_ARUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RVALID_from_SystemVerilog(  );
            axi_set_RVALID_from_SystemVerilog( _interface_ref, RVALID); // DPI call to imported task
        
        axi_propagate_RVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RVALID or posedge _check_t0_values )
    begin
        axi_local_set_RVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RLAST_from_SystemVerilog(  );
            axi_set_RLAST_from_SystemVerilog( _interface_ref, RLAST); // DPI call to imported task
        
        axi_propagate_RLAST_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RLAST or posedge _check_t0_values )
    begin
        axi_local_set_RLAST_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RDATA_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_RDATA_WIDTH ); _this_dot_1++)
        begin
            axi_set_RDATA_from_SystemVerilog_index1( _interface_ref, _this_dot_1,RDATA[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_RDATA_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RDATA or posedge _check_t0_values )
    begin
        axi_local_set_RDATA_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RRESP_from_SystemVerilog(  );
            axi_set_RRESP_from_SystemVerilog( _interface_ref, RRESP); // DPI call to imported task
        
        axi_propagate_RRESP_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RRESP or posedge _check_t0_values )
    begin
        axi_local_set_RRESP_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_RID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,RID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_RID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RID or posedge _check_t0_values )
    begin
        axi_local_set_RID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RREADY_from_SystemVerilog(  );
            axi_set_RREADY_from_SystemVerilog( _interface_ref, RREADY); // DPI call to imported task
        
        axi_propagate_RREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RREADY or posedge _check_t0_values )
    begin
        axi_local_set_RREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_RUSER_from_SystemVerilog(  );
            axi_set_RUSER_from_SystemVerilog( _interface_ref, RUSER); // DPI call to imported task
        
        axi_propagate_RUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( RUSER or posedge _check_t0_values )
    begin
        axi_local_set_RUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WVALID_from_SystemVerilog(  );
            axi_set_WVALID_from_SystemVerilog( _interface_ref, WVALID); // DPI call to imported task
        
        axi_propagate_WVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WVALID or posedge _check_t0_values )
    begin
        axi_local_set_WVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WLAST_from_SystemVerilog(  );
            axi_set_WLAST_from_SystemVerilog( _interface_ref, WLAST); // DPI call to imported task
        
        axi_propagate_WLAST_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WLAST or posedge _check_t0_values )
    begin
        axi_local_set_WLAST_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WDATA_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_WDATA_WIDTH ); _this_dot_1++)
        begin
            axi_set_WDATA_from_SystemVerilog_index1( _interface_ref, _this_dot_1,WDATA[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_WDATA_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WDATA or posedge _check_t0_values )
    begin
        axi_local_set_WDATA_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WSTRB_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( (AXI_WDATA_WIDTH / 8) ); _this_dot_1++)
        begin
            axi_set_WSTRB_from_SystemVerilog_index1( _interface_ref, _this_dot_1,WSTRB[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_WSTRB_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WSTRB or posedge _check_t0_values )
    begin
        axi_local_set_WSTRB_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_WID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,WID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_WID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WID or posedge _check_t0_values )
    begin
        axi_local_set_WID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WREADY_from_SystemVerilog(  );
            axi_set_WREADY_from_SystemVerilog( _interface_ref, WREADY); // DPI call to imported task
        
        axi_propagate_WREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WREADY or posedge _check_t0_values )
    begin
        axi_local_set_WREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_WUSER_from_SystemVerilog(  );
            axi_set_WUSER_from_SystemVerilog( _interface_ref, WUSER); // DPI call to imported task
        
        axi_propagate_WUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( WUSER or posedge _check_t0_values )
    begin
        axi_local_set_WUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BVALID_from_SystemVerilog(  );
            axi_set_BVALID_from_SystemVerilog( _interface_ref, BVALID); // DPI call to imported task
        
        axi_propagate_BVALID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BVALID or posedge _check_t0_values )
    begin
        axi_local_set_BVALID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BRESP_from_SystemVerilog(  );
            axi_set_BRESP_from_SystemVerilog( _interface_ref, BRESP); // DPI call to imported task
        
        axi_propagate_BRESP_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BRESP or posedge _check_t0_values )
    begin
        axi_local_set_BRESP_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BID_from_SystemVerilog(  );
        begin
        for (int _this_dot_1= 0; _this_dot_1 < ( AXI_ID_WIDTH ); _this_dot_1++)
        begin
            axi_set_BID_from_SystemVerilog_index1( _interface_ref, _this_dot_1,BID[_this_dot_1]); // DPI call to imported task
        
        end
        end/* 1 */ 
        axi_propagate_BID_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BID or posedge _check_t0_values )
    begin
        axi_local_set_BID_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BREADY_from_SystemVerilog(  );
            axi_set_BREADY_from_SystemVerilog( _interface_ref, BREADY); // DPI call to imported task
        
        axi_propagate_BREADY_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BREADY or posedge _check_t0_values )
    begin
        axi_local_set_BREADY_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end

    function automatic void axi_local_set_BUSER_from_SystemVerilog(  );
            axi_set_BUSER_from_SystemVerilog( _interface_ref, BUSER); // DPI call to imported task
        
        axi_propagate_BUSER_from_SystemVerilog( _interface_ref); // DPI call to imported task
    endfunction

    always @( BUSER or posedge _check_t0_values )
    begin
        axi_local_set_BUSER_from_SystemVerilog(); // Call to local task which flattens data as necessary
    end


    // CY wire and variable changed flag monitors

    always @(posedge ACLK_changed or posedge _check_t0_values )
    begin
        while (ACLK_changed == 1'b1)
        begin
            axi_get_ACLK_into_SystemVerilog( _interface_ref, internal_ACLK ); // DPI call to imported task
            ACLK_changed = 1'b0;
            #0  #0 if ( ACLK !== internal_ACLK )
            begin
                axi_local_set_ACLK_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARESETn_changed or posedge _check_t0_values )
    begin
        while (ARESETn_changed == 1'b1)
        begin
            axi_get_ARESETn_into_SystemVerilog( _interface_ref, internal_ARESETn ); // DPI call to imported task
            ARESETn_changed = 1'b0;
            #0  #0 if ( ARESETn !== internal_ARESETn )
            begin
                axi_local_set_ARESETn_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWVALID_changed or posedge _check_t0_values )
    begin
        while (AWVALID_changed == 1'b1)
        begin
            axi_get_AWVALID_into_SystemVerilog( _interface_ref, internal_AWVALID ); // DPI call to imported task
            AWVALID_changed = 1'b0;
            #0  #0 if ( AWVALID !== internal_AWVALID )
            begin
                axi_local_set_AWVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWADDR_changed or posedge _check_t0_values )
    begin
        while (AWADDR_changed == 1'b1)
        begin
            axi_get_AWADDR_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            AWADDR_changed = 1'b0;
            #0  #0 if ( AWADDR !== internal_AWADDR )
            begin
                axi_local_set_AWADDR_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWLEN_changed or posedge _check_t0_values )
    begin
        while (AWLEN_changed == 1'b1)
        begin
            axi_get_AWLEN_into_SystemVerilog( _interface_ref, internal_AWLEN ); // DPI call to imported task
            AWLEN_changed = 1'b0;
            #0  #0 if ( AWLEN !== internal_AWLEN )
            begin
                axi_local_set_AWLEN_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWSIZE_changed or posedge _check_t0_values )
    begin
        while (AWSIZE_changed == 1'b1)
        begin
            axi_get_AWSIZE_into_SystemVerilog( _interface_ref, internal_AWSIZE ); // DPI call to imported task
            AWSIZE_changed = 1'b0;
            #0  #0 if ( AWSIZE !== internal_AWSIZE )
            begin
                axi_local_set_AWSIZE_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWBURST_changed or posedge _check_t0_values )
    begin
        while (AWBURST_changed == 1'b1)
        begin
            axi_get_AWBURST_into_SystemVerilog( _interface_ref, internal_AWBURST ); // DPI call to imported task
            AWBURST_changed = 1'b0;
            #0  #0 if ( AWBURST !== internal_AWBURST )
            begin
                axi_local_set_AWBURST_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWLOCK_changed or posedge _check_t0_values )
    begin
        while (AWLOCK_changed == 1'b1)
        begin
            axi_get_AWLOCK_into_SystemVerilog( _interface_ref, internal_AWLOCK ); // DPI call to imported task
            AWLOCK_changed = 1'b0;
            #0  #0 if ( AWLOCK !== internal_AWLOCK )
            begin
                axi_local_set_AWLOCK_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWCACHE_changed or posedge _check_t0_values )
    begin
        while (AWCACHE_changed == 1'b1)
        begin
            axi_get_AWCACHE_into_SystemVerilog( _interface_ref, internal_AWCACHE ); // DPI call to imported task
            AWCACHE_changed = 1'b0;
            #0  #0 if ( AWCACHE !== internal_AWCACHE )
            begin
                axi_local_set_AWCACHE_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWPROT_changed or posedge _check_t0_values )
    begin
        while (AWPROT_changed == 1'b1)
        begin
            axi_get_AWPROT_into_SystemVerilog( _interface_ref, internal_AWPROT ); // DPI call to imported task
            AWPROT_changed = 1'b0;
            #0  #0 if ( AWPROT !== internal_AWPROT )
            begin
                axi_local_set_AWPROT_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWID_changed or posedge _check_t0_values )
    begin
        while (AWID_changed == 1'b1)
        begin
            axi_get_AWID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            AWID_changed = 1'b0;
            #0  #0 if ( AWID !== internal_AWID )
            begin
                axi_local_set_AWID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWREADY_changed or posedge _check_t0_values )
    begin
        while (AWREADY_changed == 1'b1)
        begin
            axi_get_AWREADY_into_SystemVerilog( _interface_ref, internal_AWREADY ); // DPI call to imported task
            AWREADY_changed = 1'b0;
            #0  #0 if ( AWREADY !== internal_AWREADY )
            begin
                axi_local_set_AWREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge AWUSER_changed or posedge _check_t0_values )
    begin
        while (AWUSER_changed == 1'b1)
        begin
            axi_get_AWUSER_into_SystemVerilog( _interface_ref, internal_AWUSER ); // DPI call to imported task
            AWUSER_changed = 1'b0;
            #0  #0 if ( AWUSER !== internal_AWUSER )
            begin
                axi_local_set_AWUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARVALID_changed or posedge _check_t0_values )
    begin
        while (ARVALID_changed == 1'b1)
        begin
            axi_get_ARVALID_into_SystemVerilog( _interface_ref, internal_ARVALID ); // DPI call to imported task
            ARVALID_changed = 1'b0;
            #0  #0 if ( ARVALID !== internal_ARVALID )
            begin
                axi_local_set_ARVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARADDR_changed or posedge _check_t0_values )
    begin
        while (ARADDR_changed == 1'b1)
        begin
            axi_get_ARADDR_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            ARADDR_changed = 1'b0;
            #0  #0 if ( ARADDR !== internal_ARADDR )
            begin
                axi_local_set_ARADDR_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARLEN_changed or posedge _check_t0_values )
    begin
        while (ARLEN_changed == 1'b1)
        begin
            axi_get_ARLEN_into_SystemVerilog( _interface_ref, internal_ARLEN ); // DPI call to imported task
            ARLEN_changed = 1'b0;
            #0  #0 if ( ARLEN !== internal_ARLEN )
            begin
                axi_local_set_ARLEN_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARSIZE_changed or posedge _check_t0_values )
    begin
        while (ARSIZE_changed == 1'b1)
        begin
            axi_get_ARSIZE_into_SystemVerilog( _interface_ref, internal_ARSIZE ); // DPI call to imported task
            ARSIZE_changed = 1'b0;
            #0  #0 if ( ARSIZE !== internal_ARSIZE )
            begin
                axi_local_set_ARSIZE_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARBURST_changed or posedge _check_t0_values )
    begin
        while (ARBURST_changed == 1'b1)
        begin
            axi_get_ARBURST_into_SystemVerilog( _interface_ref, internal_ARBURST ); // DPI call to imported task
            ARBURST_changed = 1'b0;
            #0  #0 if ( ARBURST !== internal_ARBURST )
            begin
                axi_local_set_ARBURST_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARLOCK_changed or posedge _check_t0_values )
    begin
        while (ARLOCK_changed == 1'b1)
        begin
            axi_get_ARLOCK_into_SystemVerilog( _interface_ref, internal_ARLOCK ); // DPI call to imported task
            ARLOCK_changed = 1'b0;
            #0  #0 if ( ARLOCK !== internal_ARLOCK )
            begin
                axi_local_set_ARLOCK_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARCACHE_changed or posedge _check_t0_values )
    begin
        while (ARCACHE_changed == 1'b1)
        begin
            axi_get_ARCACHE_into_SystemVerilog( _interface_ref, internal_ARCACHE ); // DPI call to imported task
            ARCACHE_changed = 1'b0;
            #0  #0 if ( ARCACHE !== internal_ARCACHE )
            begin
                axi_local_set_ARCACHE_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARPROT_changed or posedge _check_t0_values )
    begin
        while (ARPROT_changed == 1'b1)
        begin
            axi_get_ARPROT_into_SystemVerilog( _interface_ref, internal_ARPROT ); // DPI call to imported task
            ARPROT_changed = 1'b0;
            #0  #0 if ( ARPROT !== internal_ARPROT )
            begin
                axi_local_set_ARPROT_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARID_changed or posedge _check_t0_values )
    begin
        while (ARID_changed == 1'b1)
        begin
            axi_get_ARID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            ARID_changed = 1'b0;
            #0  #0 if ( ARID !== internal_ARID )
            begin
                axi_local_set_ARID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARREADY_changed or posedge _check_t0_values )
    begin
        while (ARREADY_changed == 1'b1)
        begin
            axi_get_ARREADY_into_SystemVerilog( _interface_ref, internal_ARREADY ); // DPI call to imported task
            ARREADY_changed = 1'b0;
            #0  #0 if ( ARREADY !== internal_ARREADY )
            begin
                axi_local_set_ARREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge ARUSER_changed or posedge _check_t0_values )
    begin
        while (ARUSER_changed == 1'b1)
        begin
            axi_get_ARUSER_into_SystemVerilog( _interface_ref, internal_ARUSER ); // DPI call to imported task
            ARUSER_changed = 1'b0;
            #0  #0 if ( ARUSER !== internal_ARUSER )
            begin
                axi_local_set_ARUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RVALID_changed or posedge _check_t0_values )
    begin
        while (RVALID_changed == 1'b1)
        begin
            axi_get_RVALID_into_SystemVerilog( _interface_ref, internal_RVALID ); // DPI call to imported task
            RVALID_changed = 1'b0;
            #0  #0 if ( RVALID !== internal_RVALID )
            begin
                axi_local_set_RVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RLAST_changed or posedge _check_t0_values )
    begin
        while (RLAST_changed == 1'b1)
        begin
            axi_get_RLAST_into_SystemVerilog( _interface_ref, internal_RLAST ); // DPI call to imported task
            RLAST_changed = 1'b0;
            #0  #0 if ( RLAST !== internal_RLAST )
            begin
                axi_local_set_RLAST_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RDATA_changed or posedge _check_t0_values )
    begin
        while (RDATA_changed == 1'b1)
        begin
            axi_get_RDATA_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            RDATA_changed = 1'b0;
            #0  #0 if ( RDATA !== internal_RDATA )
            begin
                axi_local_set_RDATA_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RRESP_changed or posedge _check_t0_values )
    begin
        while (RRESP_changed == 1'b1)
        begin
            axi_get_RRESP_into_SystemVerilog( _interface_ref, internal_RRESP ); // DPI call to imported task
            RRESP_changed = 1'b0;
            #0  #0 if ( RRESP !== internal_RRESP )
            begin
                axi_local_set_RRESP_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RID_changed or posedge _check_t0_values )
    begin
        while (RID_changed == 1'b1)
        begin
            axi_get_RID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            RID_changed = 1'b0;
            #0  #0 if ( RID !== internal_RID )
            begin
                axi_local_set_RID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RREADY_changed or posedge _check_t0_values )
    begin
        while (RREADY_changed == 1'b1)
        begin
            axi_get_RREADY_into_SystemVerilog( _interface_ref, internal_RREADY ); // DPI call to imported task
            RREADY_changed = 1'b0;
            #0  #0 if ( RREADY !== internal_RREADY )
            begin
                axi_local_set_RREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge RUSER_changed or posedge _check_t0_values )
    begin
        while (RUSER_changed == 1'b1)
        begin
            axi_get_RUSER_into_SystemVerilog( _interface_ref, internal_RUSER ); // DPI call to imported task
            RUSER_changed = 1'b0;
            #0  #0 if ( RUSER !== internal_RUSER )
            begin
                axi_local_set_RUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WVALID_changed or posedge _check_t0_values )
    begin
        while (WVALID_changed == 1'b1)
        begin
            axi_get_WVALID_into_SystemVerilog( _interface_ref, internal_WVALID ); // DPI call to imported task
            WVALID_changed = 1'b0;
            #0  #0 if ( WVALID !== internal_WVALID )
            begin
                axi_local_set_WVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WLAST_changed or posedge _check_t0_values )
    begin
        while (WLAST_changed == 1'b1)
        begin
            axi_get_WLAST_into_SystemVerilog( _interface_ref, internal_WLAST ); // DPI call to imported task
            WLAST_changed = 1'b0;
            #0  #0 if ( WLAST !== internal_WLAST )
            begin
                axi_local_set_WLAST_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WDATA_changed or posedge _check_t0_values )
    begin
        while (WDATA_changed == 1'b1)
        begin
            axi_get_WDATA_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            WDATA_changed = 1'b0;
            #0  #0 if ( WDATA !== internal_WDATA )
            begin
                axi_local_set_WDATA_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WSTRB_changed or posedge _check_t0_values )
    begin
        while (WSTRB_changed == 1'b1)
        begin
            axi_get_WSTRB_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            WSTRB_changed = 1'b0;
            #0  #0 if ( WSTRB !== internal_WSTRB )
            begin
                axi_local_set_WSTRB_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WID_changed or posedge _check_t0_values )
    begin
        while (WID_changed == 1'b1)
        begin
            axi_get_WID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            WID_changed = 1'b0;
            #0  #0 if ( WID !== internal_WID )
            begin
                axi_local_set_WID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WREADY_changed or posedge _check_t0_values )
    begin
        while (WREADY_changed == 1'b1)
        begin
            axi_get_WREADY_into_SystemVerilog( _interface_ref, internal_WREADY ); // DPI call to imported task
            WREADY_changed = 1'b0;
            #0  #0 if ( WREADY !== internal_WREADY )
            begin
                axi_local_set_WREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge WUSER_changed or posedge _check_t0_values )
    begin
        while (WUSER_changed == 1'b1)
        begin
            axi_get_WUSER_into_SystemVerilog( _interface_ref, internal_WUSER ); // DPI call to imported task
            WUSER_changed = 1'b0;
            #0  #0 if ( WUSER !== internal_WUSER )
            begin
                axi_local_set_WUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BVALID_changed or posedge _check_t0_values )
    begin
        while (BVALID_changed == 1'b1)
        begin
            axi_get_BVALID_into_SystemVerilog( _interface_ref, internal_BVALID ); // DPI call to imported task
            BVALID_changed = 1'b0;
            #0  #0 if ( BVALID !== internal_BVALID )
            begin
                axi_local_set_BVALID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BRESP_changed or posedge _check_t0_values )
    begin
        while (BRESP_changed == 1'b1)
        begin
            axi_get_BRESP_into_SystemVerilog( _interface_ref, internal_BRESP ); // DPI call to imported task
            BRESP_changed = 1'b0;
            #0  #0 if ( BRESP !== internal_BRESP )
            begin
                axi_local_set_BRESP_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BID_changed or posedge _check_t0_values )
    begin
        while (BID_changed == 1'b1)
        begin
            axi_get_BID_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            BID_changed = 1'b0;
            #0  #0 if ( BID !== internal_BID )
            begin
                axi_local_set_BID_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BREADY_changed or posedge _check_t0_values )
    begin
        while (BREADY_changed == 1'b1)
        begin
            axi_get_BREADY_into_SystemVerilog( _interface_ref, internal_BREADY ); // DPI call to imported task
            BREADY_changed = 1'b0;
            #0  #0 if ( BREADY !== internal_BREADY )
            begin
                axi_local_set_BREADY_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge BUSER_changed or posedge _check_t0_values )
    begin
        while (BUSER_changed == 1'b1)
        begin
            axi_get_BUSER_into_SystemVerilog( _interface_ref, internal_BUSER ); // DPI call to imported task
            BUSER_changed = 1'b0;
            #0  #0 if ( BUSER !== internal_BUSER )
            begin
                axi_local_set_BUSER_from_SystemVerilog(  );
            end
        end
    end

    always @(posedge config_write_ctrl_to_data_mintime_changed or posedge _check_t0_values )
    begin
        if (config_write_ctrl_to_data_mintime_changed == 1'b1)
        begin
            axi_get_config_write_ctrl_to_data_mintime_into_SystemVerilog( _interface_ref, config_write_ctrl_to_data_mintime ); // DPI call to imported task
            config_write_ctrl_to_data_mintime_changed = 1'b0;
        end
    end

    always @(posedge config_master_write_delay_changed or posedge _check_t0_values )
    begin
        if (config_master_write_delay_changed == 1'b1)
        begin
            axi_get_config_master_write_delay_into_SystemVerilog( _interface_ref, config_master_write_delay ); // DPI call to imported task
            config_master_write_delay_changed = 1'b0;
        end
    end

    always @(posedge config_enable_all_assertions_changed or posedge _check_t0_values )
    begin
        if (config_enable_all_assertions_changed == 1'b1)
        begin
            axi_get_config_enable_all_assertions_into_SystemVerilog( _interface_ref, config_enable_all_assertions ); // DPI call to imported task
            config_enable_all_assertions_changed = 1'b0;
        end
    end

    always @(posedge config_enable_assertion_changed or posedge _check_t0_values )
    begin
        if (config_enable_assertion_changed == 1'b1)
        begin
            axi_get_config_enable_assertion_into_SystemVerilog( _interface_ref, config_enable_assertion ); // DPI call to imported task
            config_enable_assertion_changed = 1'b0;
        end
    end

    always @(posedge config_slave_start_addr_changed or posedge _check_t0_values )
    begin
        if (config_slave_start_addr_changed == 1'b1)
        begin
            axi_get_config_slave_start_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            config_slave_start_addr_changed = 1'b0;
        end
    end

    always @(posedge config_slave_end_addr_changed or posedge _check_t0_values )
    begin
        if (config_slave_end_addr_changed == 1'b1)
        begin
            axi_get_config_slave_end_addr_into_SystemVerilog( _interface_ref ); // DPI call to imported task
            config_slave_end_addr_changed = 1'b0;
        end
    end

    always @(posedge config_support_exclusive_access_changed or posedge _check_t0_values )
    begin
        if (config_support_exclusive_access_changed == 1'b1)
        begin
            axi_get_config_support_exclusive_access_into_SystemVerilog( _interface_ref, config_support_exclusive_access ); // DPI call to imported task
            config_support_exclusive_access_changed = 1'b0;
        end
    end

    always @(posedge config_read_data_reordering_depth_changed or posedge _check_t0_values )
    begin
        if (config_read_data_reordering_depth_changed == 1'b1)
        begin
            axi_get_config_read_data_reordering_depth_into_SystemVerilog( _interface_ref, config_read_data_reordering_depth ); // DPI call to imported task
            config_read_data_reordering_depth_changed = 1'b0;
        end
    end

    always @(posedge config_max_transaction_time_factor_changed or posedge _check_t0_values )
    begin
        if (config_max_transaction_time_factor_changed == 1'b1)
        begin
            axi_get_config_max_transaction_time_factor_into_SystemVerilog( _interface_ref, config_max_transaction_time_factor ); // DPI call to imported task
            config_max_transaction_time_factor_changed = 1'b0;
        end
    end

    always @(posedge config_timeout_max_data_transfer_changed or posedge _check_t0_values )
    begin
        if (config_timeout_max_data_transfer_changed == 1'b1)
        begin
            axi_get_config_timeout_max_data_transfer_into_SystemVerilog( _interface_ref, config_timeout_max_data_transfer ); // DPI call to imported task
            config_timeout_max_data_transfer_changed = 1'b0;
        end
    end

    always @(posedge config_burst_timeout_factor_changed or posedge _check_t0_values )
    begin
        if (config_burst_timeout_factor_changed == 1'b1)
        begin
            axi_get_config_burst_timeout_factor_into_SystemVerilog( _interface_ref, config_burst_timeout_factor ); // DPI call to imported task
            config_burst_timeout_factor_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_AWVALID_assertion_to_AWREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_AWVALID_assertion_to_AWREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_AWVALID_assertion_to_AWREADY_into_SystemVerilog( _interface_ref, config_max_latency_AWVALID_assertion_to_AWREADY ); // DPI call to imported task
            config_max_latency_AWVALID_assertion_to_AWREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_ARVALID_assertion_to_ARREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_ARVALID_assertion_to_ARREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_ARVALID_assertion_to_ARREADY_into_SystemVerilog( _interface_ref, config_max_latency_ARVALID_assertion_to_ARREADY ); // DPI call to imported task
            config_max_latency_ARVALID_assertion_to_ARREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_RVALID_assertion_to_RREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_RVALID_assertion_to_RREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_RVALID_assertion_to_RREADY_into_SystemVerilog( _interface_ref, config_max_latency_RVALID_assertion_to_RREADY ); // DPI call to imported task
            config_max_latency_RVALID_assertion_to_RREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_BVALID_assertion_to_BREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_BVALID_assertion_to_BREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_BVALID_assertion_to_BREADY_into_SystemVerilog( _interface_ref, config_max_latency_BVALID_assertion_to_BREADY ); // DPI call to imported task
            config_max_latency_BVALID_assertion_to_BREADY_changed = 1'b0;
        end
    end

    always @(posedge config_max_latency_WVALID_assertion_to_WREADY_changed or posedge _check_t0_values )
    begin
        if (config_max_latency_WVALID_assertion_to_WREADY_changed == 1'b1)
        begin
            axi_get_config_max_latency_WVALID_assertion_to_WREADY_into_SystemVerilog( _interface_ref, config_max_latency_WVALID_assertion_to_WREADY ); // DPI call to imported task
            config_max_latency_WVALID_assertion_to_WREADY_changed = 1'b0;
        end
    end

    always @(posedge config_master_error_position_changed or posedge _check_t0_values )
    begin
        if (config_master_error_position_changed == 1'b1)
        begin
            axi_get_config_master_error_position_into_SystemVerilog( _interface_ref, config_master_error_position ); // DPI call to imported task
            config_master_error_position_changed = 1'b0;
        end
    end

    always @(posedge config_setup_time_changed or posedge _check_t0_values )
    begin
        if (config_setup_time_changed == 1'b1)
        begin
            axi_get_config_setup_time_into_SystemVerilog( _interface_ref, config_setup_time ); // DPI call to imported task
            config_setup_time_changed = 1'b0;
        end
    end

    always @(posedge config_hold_time_changed or posedge _check_t0_values )
    begin
        if (config_hold_time_changed == 1'b1)
        begin
            axi_get_config_hold_time_into_SystemVerilog( _interface_ref, config_hold_time ); // DPI call to imported task
            config_hold_time_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_wr_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_wr_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_wr_into_SystemVerilog( _interface_ref, config_max_outstanding_wr ); // DPI call to imported task
            config_max_outstanding_wr_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_rd_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_rd_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_rd_into_SystemVerilog( _interface_ref, config_max_outstanding_rd ); // DPI call to imported task
            config_max_outstanding_rd_changed = 1'b0;
        end
    end

    always @(posedge config_max_outstanding_rw_changed or posedge _check_t0_values )
    begin
        if (config_max_outstanding_rw_changed == 1'b1)
        begin
            axi_get_config_max_outstanding_rw_into_SystemVerilog( _interface_ref, config_max_outstanding_rw ); // DPI call to imported task
            config_max_outstanding_rw_changed = 1'b0;
        end
    end

    always @(posedge config_is_issuing_changed or posedge _check_t0_values )
    begin
        if (config_is_issuing_changed == 1'b1)
        begin
            axi_get_config_is_issuing_into_SystemVerilog( _interface_ref, config_is_issuing ); // DPI call to imported task
            config_is_issuing_changed = 1'b0;
        end
    end


    //--------------------------------------------------------------------------------
    // Task which blocks and outputs an error if the interface has not initialized properly
    //--------------------------------------------------------------------------------

    task _initialized();
        if (_interface_ref == 0)
        begin
            $display("Error: %m - Questa Verification IP failed to initialise. Please check questa_mvc.log for details");
            wait(_interface_ref!=0);
        end
    endtask

endinterface

`endif // VCS
