module interrupt_handler(
    input clk, rst,
    input external,
    output [31:0] interrupt_handling_addr,
    output interrupt_ctrl
);
    
endmodule